module systemcdes (
x1710,
x1826,
x1244,
x815,
x761,
x2017,
x1785,
x843,
x1024,
x2211,
x997,
x1361,
x748,
x1800,
x1636,
x876,
x1742,
x621,
x1517,
x1435,
x1681,
x597,
x3333,
x1262,
x523,
x1490,
x1007,
x780,
x42206,
x1662,
x2480,
x1427,
x497,
x1286,
x717,
x692,
x850,
x1186,
x585,
x1456,
x1318,
x1844,
x535,
x42204,
x1808,
x554,
x651,
x1466,
x1980,
x808,
x1047,
x914,
x1750,
x945,
x857,
x972,
x629,
x1645,
x1086,
x2269,
x2143,
x831,
x562,
x675,
x793,
x935,
x1582,
x1110,
x1593,
x663,
x1958,
x1889,
x1031,
x1192,
x956,
x1546,
x42209,
x1063,
x899,
x1719,
x1611,
x921,
x42207,
x990,
x2242,
x883,
x1312,
x1280,
x1877,
x42202,
x1554,
x515,
x2062,
x2167,
x543,
x1915,
x1343,
x2116,
x730,
x1126,
x506,
x1170,
x1835,
x1368,
x1868,
x2080,
x2183,
x1620,
x1769,
x609,
x1933,
x42203,
x638,
x1863,
x2026,
x2049,
x1381,
x42208,
x1993,
x1014,
x1073,
x870,
x701,
x1214,
x1146,
x1222,
x1817,
x574,
x1405,
x1333,
x1851,
x42205,
x397,
x363,
x279,
x237,
x451,
x266,
x444,
x355,
x185,
x439,
x429,
x44,
x128,
x378,
x216,
x177,
x193,
x316,
x152,
x459,
x467,
x64,
x90,
x201,
x347,
x245,
x114,
x144,
x309,
x331,
x136,
x170,
x405,
x10,
x72,
x121,
x339,
x434,
x229,
x302,
x370,
x20,
x98,
x223,
x295,
x421,
x31,
x0,
x258,
x413,
x166,
x57,
x106,
x36,
x484,
x208,
x78,
x49,
x273,
x389,
x323,
x83,
x253,
x287,
x159);

// Start PIs
input x1710;
input x1826;
input x1244;
input x815;
input x761;
input x2017;
input x1785;
input x843;
input x1024;
input x2211;
input x997;
input x1361;
input x748;
input x1800;
input x1636;
input x876;
input x1742;
input x621;
input x1517;
input x1435;
input x1681;
input x597;
input x3333;
input x1262;
input x523;
input x1490;
input x1007;
input x780;
input x42206;
input x1662;
input x2480;
input x1427;
input x497;
input x1286;
input x717;
input x692;
input x850;
input x1186;
input x585;
input x1456;
input x1318;
input x1844;
input x535;
input x42204;
input x1808;
input x554;
input x651;
input x1466;
input x1980;
input x808;
input x1047;
input x914;
input x1750;
input x945;
input x857;
input x972;
input x629;
input x1645;
input x1086;
input x2269;
input x2143;
input x831;
input x562;
input x675;
input x793;
input x935;
input x1582;
input x1110;
input x1593;
input x663;
input x1958;
input x1889;
input x1031;
input x1192;
input x956;
input x1546;
input x42209;
input x1063;
input x899;
input x1719;
input x1611;
input x921;
input x42207;
input x990;
input x2242;
input x883;
input x1312;
input x1280;
input x1877;
input x42202;
input x1554;
input x515;
input x2062;
input x2167;
input x543;
input x1915;
input x1343;
input x2116;
input x730;
input x1126;
input x506;
input x1170;
input x1835;
input x1368;
input x1868;
input x2080;
input x2183;
input x1620;
input x1769;
input x609;
input x1933;
input x42203;
input x638;
input x1863;
input x2026;
input x2049;
input x1381;
input x42208;
input x1993;
input x1014;
input x1073;
input x870;
input x701;
input x1214;
input x1146;
input x1222;
input x1817;
input x574;
input x1405;
input x1333;
input x1851;
input x42205;

// Start POs
output x397;
output x363;
output x279;
output x237;
output x451;
output x266;
output x444;
output x355;
output x185;
output x439;
output x429;
output x44;
output x128;
output x378;
output x216;
output x177;
output x193;
output x316;
output x152;
output x459;
output x467;
output x64;
output x90;
output x201;
output x347;
output x245;
output x114;
output x144;
output x309;
output x331;
output x136;
output x170;
output x405;
output x10;
output x72;
output x121;
output x339;
output x434;
output x229;
output x302;
output x370;
output x20;
output x98;
output x223;
output x295;
output x421;
output x31;
output x0;
output x258;
output x413;
output x166;
output x57;
output x106;
output x36;
output x484;
output x208;
output x78;
output x49;
output x273;
output x389;
output x323;
output x83;
output x253;
output x287;
output x159;

// Start wires
wire net_2388;
wire net_2449;
wire net_1317;
wire net_416;
wire net_215;
wire net_2394;
wire net_933;
wire net_2418;
wire net_1382;
wire net_1244;
wire net_1215;
wire net_943;
wire net_429;
wire net_3377;
wire net_129;
wire net_373;
wire net_98;
wire net_1897;
wire net_980;
wire net_151;
wire net_356;
wire net_53;
wire net_2542;
wire x843;
wire net_1786;
wire net_1377;
wire net_1625;
wire net_452;
wire x1024;
wire x2211;
wire net_545;
wire net_2147;
wire net_1483;
wire net_284;
wire net_560;
wire net_3031;
wire net_439;
wire net_2513;
wire net_259;
wire net_3351;
wire net_2645;
wire net_1393;
wire net_2169;
wire net_3119;
wire net_1324;
wire net_1231;
wire net_187;
wire net_2256;
wire x1435;
wire x3333;
wire net_264;
wire net_3305;
wire net_2207;
wire net_2674;
wire net_263;
wire net_2872;
wire net_1138;
wire net_160;
wire net_2432;
wire net_2769;
wire net_832;
wire net_322;
wire net_1671;
wire net_1064;
wire net_815;
wire net_2082;
wire net_420;
wire net_3292;
wire net_1746;
wire net_1439;
wire net_665;
wire x170;
wire net_2222;
wire x717;
wire net_1778;
wire net_508;
wire net_2825;
wire net_2322;
wire net_1090;
wire net_586;
wire net_1347;
wire net_1091;
wire net_3341;
wire net_703;
wire net_1072;
wire net_193;
wire net_120;
wire net_292;
wire net_201;
wire net_1706;
wire net_109;
wire net_2942;
wire net_3280;
wire net_3085;
wire net_96;
wire net_1730;
wire net_2921;
wire net_2896;
wire net_3281;
wire net_167;
wire net_3289;
wire net_651;
wire net_3134;
wire net_2931;
wire net_1852;
wire net_3415;
wire net_3114;
wire net_1720;
wire net_744;
wire net_2556;
wire net_1555;
wire net_598;
wire net_2060;
wire net_2051;
wire net_2780;
wire net_2740;
wire net_789;
wire x323;
wire net_2806;
wire net_2011;
wire net_3244;
wire net_593;
wire net_672;
wire net_2171;
wire net_777;
wire net_2765;
wire net_3157;
wire net_2820;
wire net_2027;
wire net_490;
wire net_742;
wire x266;
wire net_3068;
wire net_2425;
wire net_2456;
wire net_2753;
wire net_2830;
wire net_1232;
wire net_1198;
wire net_2509;
wire net_1953;
wire net_3059;
wire net_2862;
wire net_1860;
wire net_632;
wire net_2457;
wire net_883;
wire net_843;
wire net_2156;
wire net_1432;
wire net_464;
wire net_2841;
wire net_1312;
wire net_2957;
wire net_1977;
wire net_446;
wire net_2100;
wire net_2938;
wire net_2122;
wire net_1516;
wire net_1712;
wire net_1171;
wire net_1540;
wire net_248;
wire net_3063;
wire net_1083;
wire net_3343;
wire x309;
wire net_3423;
wire net_1499;
wire net_964;
wire net_3326;
wire net_1453;
wire net_2913;
wire net_1725;
wire net_3295;
wire net_2239;
wire net_3394;
wire net_2268;
wire net_1256;
wire net_634;
wire net_1413;
wire net_802;
wire x339;
wire x1620;
wire net_2846;
wire net_2303;
wire net_371;
wire net_1735;
wire net_2787;
wire net_1767;
wire net_3041;
wire net_2210;
wire net_1840;
wire net_2176;
wire net_1571;
wire net_1640;
wire x2026;
wire net_2466;
wire net_2724;
wire net_997;
wire net_1031;
wire net_1741;
wire net_503;
wire net_256;
wire net_850;
wire net_1140;
wire net_2764;
wire net_2103;
wire net_1672;
wire net_1636;
wire net_1464;
wire net_996;
wire net_3257;
wire net_3091;
wire net_679;
wire net_2994;
wire net_1168;
wire net_2680;
wire net_3196;
wire net_308;
wire net_75;
wire net_959;
wire net_515;
wire net_1334;
wire net_757;
wire net_206;
wire net_3051;
wire net_2020;
wire net_1688;
wire net_3090;
wire net_2345;
wire net_223;
wire net_1009;
wire net_715;
wire net_235;
wire net_2973;
wire net_2077;
wire net_890;
wire net_3106;
wire net_2219;
wire net_2745;
wire net_2546;
wire net_2961;
wire net_2503;
wire net_2374;
wire net_2164;
wire net_1876;
wire net_2471;
wire net_250;
wire net_3081;
wire net_312;
wire net_2404;
wire net_130;
wire net_2627;
wire net_572;
wire net_2055;
wire net_147;
wire net_481;
wire net_369;
wire net_2630;
wire net_1662;
wire net_2338;
wire net_1985;
wire net_403;
wire net_2340;
wire net_2616;
wire net_1079;
wire net_32;
wire net_2444;
wire net_1596;
wire net_282;
wire net_2275;
wire net_2809;
wire net_1188;
wire net_3235;
wire net_780;
wire net_3184;
wire net_1446;
wire net_841;
wire net_541;
wire net_1750;
wire net_794;
wire net_2397;
wire net_2370;
wire net_3346;
wire net_2047;
wire net_2469;
wire net_1251;
wire net_2693;
wire net_2391;
wire net_528;
wire net_2802;
wire net_2906;
wire net_1404;
wire net_1012;
wire net_456;
wire net_155;
wire net_1697;
wire net_335;
wire net_1468;
wire net_907;
wire net_181;
wire net_1753;
wire net_3333;
wire net_349;
wire net_39;
wire net_3076;
wire net_2435;
wire net_245;
wire net_1409;
wire net_2383;
wire x370;
wire net_2036;
wire net_395;
wire net_2539;
wire net_2977;
wire net_1130;
wire net_493;
wire net_2719;
wire net_386;
wire net_2323;
wire net_1428;
wire net_987;
wire net_641;
wire net_277;
wire net_1965;
wire net_1790;
wire net_2798;
wire net_89;
wire net_1152;
wire net_3071;
wire net_2350;
wire net_2318;
wire net_1226;
wire net_3271;
wire net_680;
wire net_1901;
wire net_3021;
wire net_338;
wire net_1039;
wire net_2998;
wire net_1709;
wire net_721;
wire net_243;
wire net_3226;
wire net_3143;
wire net_400;
wire net_1935;
wire net_2757;
wire net_1018;
wire net_602;
wire net_2854;
wire net_2379;
wire net_2009;
wire net_2369;
wire net_2038;
wire net_1818;
wire net_175;
wire net_2918;
wire net_823;
wire net_2925;
wire net_1850;
wire net_1497;
wire net_106;
wire net_1800;
wire net_1380;
wire net_1676;
wire net_1855;
wire net_279;
wire net_3347;
wire net_1992;
wire net_1523;
wire net_1177;
wire net_1163;
wire net_698;
wire net_1656;
wire net_897;
wire net_1915;
wire net_1191;
wire net_2853;
wire net_2255;
wire net_691;
wire net_2705;
wire x1546;
wire net_615;
wire net_2485;
wire net_3273;
wire net_1997;
wire net_3178;
wire net_1559;
wire net_441;
wire net_2701;
wire net_2833;
wire net_1863;
wire net_1620;
wire net_2608;
wire net_138;
wire net_749;
wire net_2561;
wire net_1019;
wire net_2813;
wire net_2663;
wire net_1948;
wire net_1616;
wire net_728;
wire net_1276;
wire net_1006;
wire net_719;
wire net_2781;
wire net_2519;
wire net_170;
wire net_471;
wire net_2571;
wire net_1055;
wire net_1531;
wire net_878;
wire net_1159;
wire net_2969;
wire net_518;
wire net_861;
wire net_57;
wire net_3222;
wire net_929;
wire net_3321;
wire net_1418;
wire net_3202;
wire net_2523;
wire net_708;
wire net_2985;
wire net_696;
wire net_537;
wire net_3216;
wire net_3056;
wire net_1565;
wire net_1713;
wire net_169;
wire net_2668;
wire net_171;
wire net_2677;
wire x1381;
wire net_3252;
wire net_2775;
wire net_2234;
wire net_513;
wire net_604;
wire net_163;
wire net_967;
wire net_1576;
wire net_1421;
wire net_1527;
wire net_268;
wire net_3407;
wire net_2736;
wire net_2127;
wire net_1280;
wire net_459;
wire net_3386;
wire net_483;
wire net_48;
wire net_1149;
wire net_737;
wire net_2284;
wire net_3412;
wire net_2962;
wire net_2113;
wire net_1645;
wire net_2193;
wire net_176;
wire net_2570;
wire net_1298;
wire net_296;
wire net_2131;
wire net_3354;
wire net_614;
wire net_2712;
wire net_2005;
wire net_2771;
wire net_1886;
wire net_1156;
wire net_1123;
wire net_3194;
wire net_2604;
wire x997;
wire net_2228;
wire net_1966;
wire net_3020;
wire net_786;
wire net_1192;
wire net_127;
wire net_3363;
wire net_1339;
wire net_984;
wire net_1105;
wire net_101;
wire net_906;
wire net_1659;
wire net_1272;
wire net_3156;
wire net_2422;
wire net_2172;
wire net_326;
wire net_2482;
wire net_2381;
wire net_2109;
wire net_1770;
wire net_707;
wire net_589;
wire x90;
wire net_655;
wire x1007;
wire net_652;
wire net_1814;
wire net_1815;
wire net_1856;
wire net_830;
wire net_3175;
wire net_2505;
wire net_575;
wire net_1279;
wire net_877;
wire net_378;
wire net_2829;
wire net_1047;
wire net_724;
wire net_3309;
wire net_2799;
wire net_3142;
wire net_3036;
wire net_423;
wire net_1219;
wire net_328;
wire net_2683;
wire net_2631;
wire net_2384;
wire net_1958;
wire net_1931;
wire net_2877;
wire net_2165;
wire net_2480;
wire net_3294;
wire net_1549;
wire net_3284;
wire net_3016;
wire net_1474;
wire net_1467;
wire net_3181;
wire net_2784;
wire net_1061;
wire net_874;
wire net_2929;
wire net_1632;
wire net_765;
wire net_675;
wire net_2562;
wire net_1342;
wire net_2867;
wire net_2633;
wire net_1661;
wire net_1666;
wire net_1236;
wire net_818;
wire net_2288;
wire net_2746;
wire net_2700;
wire net_2099;
wire net_1211;
wire net_2182;
wire net_1768;
wire net_1183;
wire net_2594;
wire net_150;
wire net_1488;
wire net_2812;
wire net_304;
wire net_1684;
wire net_811;
wire net_352;
wire net_30;
wire net_2021;
wire net_1703;
wire net_1068;
wire net_1462;
wire net_436;
wire net_2837;
wire net_186;
wire net_2017;
wire net_2495;
wire net_2824;
wire net_1777;
wire net_1926;
wire net_3115;
wire net_2735;
wire net_1050;
wire net_2760;
wire net_2072;
wire net_1641;
wire net_1316;
wire x177;
wire net_1872;
wire net_2271;
wire net_1621;
wire net_792;
wire net_3070;
wire net_3409;
wire net_2203;
wire net_1904;
wire net_1716;
wire net_1702;
wire net_1103;
wire net_1035;
wire net_767;
wire net_1607;
wire net_3055;
wire net_1838;
wire net_219;
wire net_1263;
wire net_2187;
wire net_131;
wire net_2476;
wire net_196;
wire net_913;
wire net_2067;
wire net_358;
wire net_1973;
wire net_3130;
wire net_3095;
wire net_2845;
wire net_2016;
wire net_2934;
wire net_3387;
wire net_2641;
wire net_1479;
wire net_1763;
wire net_1639;
wire net_3125;
wire net_3094;
wire x1126;
wire net_1285;
wire net_360;
wire net_3112;
wire net_1927;
wire net_1175;
wire net_213;
wire net_2882;
wire net_2324;
wire net_3278;
wire net_260;
wire net_2947;
wire net_2922;
wire net_947;
wire net_3137;
wire net_1513;
wire net_2152;
wire net_1126;
wire net_732;
wire net_2004;
wire net_1742;
wire net_3064;
wire net_1325;
wire net_2276;
wire net_3316;
wire net_3032;
wire net_1597;
wire net_1373;
wire net_1352;
wire net_2885;
wire net_2567;
wire net_2088;
wire net_468;
wire x1146;
wire net_1187;
wire net_2689;
wire net_798;
wire net_3135;
wire net_2761;
wire net_73;
wire net_3206;
wire net_2059;
wire net_1303;
wire net_2858;
wire net_3370;
wire net_1899;
wire net_1503;
wire net_1336;
wire net_2102;
wire net_179;
wire net_61;
wire net_1843;
wire net_1442;
wire net_449;
wire net_1807;
wire net_62;
wire net_1943;
wire net_1930;
wire net_3261;
wire net_534;
wire net_1087;
wire net_733;
wire net_3336;
wire net_887;
wire x2017;
wire net_2289;
wire net_903;
wire net_1551;
wire net_486;
wire net_1894;
wire net_2031;
wire net_1868;
wire net_1560;
wire net_406;
wire x193;
wire net_2431;
wire net_2308;
wire net_2378;
wire net_633;
wire net_113;
wire net_2989;
wire net_497;
wire net_1914;
wire net_40;
wire net_2770;
wire net_2408;
wire net_2636;
wire net_1424;
wire net_1414;
wire net_300;
wire net_2652;
wire net_3382;
wire net_2720;
wire net_1545;
wire net_1457;
wire net_1233;
wire net_748;
wire x2480;
wire net_2741;
wire net_95;
wire net_1834;
wire net_990;
wire net_950;
wire x405;
wire net_2448;
wire net_1436;
wire net_2327;
wire net_1003;
wire net_514;
wire net_2332;
wire x72;
wire net_1604;
wire net_2715;
wire net_1803;
wire net_3400;
wire net_1941;
wire net_3392;
wire net_524;
wire net_2551;
wire net_2816;
wire net_1134;
wire net_646;
wire net_363;
wire net_2731;
wire net_445;
wire net_2601;
wire net_1319;
wire net_1214;
wire net_776;
wire net_3080;
wire net_866;
wire net_2891;
wire net_2508;
wire net_44;
wire net_1650;
wire net_1582;
wire net_520;
wire x31;
wire net_3150;
wire net_3149;
wire net_1675;
wire net_1032;
wire net_2247;
wire net_567;
wire x945;
wire net_2333;
wire net_2213;
wire net_3231;
wire net_1368;
wire net_981;
wire net_2575;
wire net_272;
wire net_1248;
wire net_2401;
wire net_2291;
wire net_1097;
wire net_2238;
wire net_845;
wire net_1024;
wire x287;
wire net_1590;
wire net_1566;
wire x1086;
wire net_762;
wire net_1305;
wire x831;
wire net_2354;
wire net_1612;
wire net_695;
wire net_839;
wire net_1387;
wire net_2525;
wire net_1201;
wire net_814;
wire net_1581;
wire net_556;
wire net_2671;
wire net_3330;
wire net_893;
wire net_2413;
wire net_559;
wire net_255;
wire net_3042;
wire net_2792;
wire net_345;
wire net_2965;
wire net_2128;
wire net_1717;
wire net_859;
wire net_620;
wire net_3299;
wire net_2586;
wire net_619;
wire net_1167;
wire net_1655;
wire net_398;
wire net_3399;
wire net_2365;
wire net_954;
wire net_2198;
wire net_1044;
wire net_2117;
wire net_2461;
wire net_1766;
wire net_2940;
wire net_2582;
wire net_2043;
wire net_2095;
wire net_2598;
wire net_2361;
wire net_3285;
wire net_2879;
wire net_1572;
wire net_1680;
wire net_68;
wire net_2314;
wire net_2613;
wire net_3302;
wire net_1493;
wire net_976;
wire net_3187;
wire net_2134;
wire net_2709;
wire net_2622;
wire x10;
wire net_316;
wire net_865;
wire net_84;
wire net_611;
wire net_231;
wire net_2621;
wire net_2579;
wire net_3024;
wire net_1223;
wire net_2750;
wire net_1759;
wire net_1866;
wire net_2262;
wire net_926;
wire net_3011;
wire net_3211;
wire net_2160;
wire net_2087;
wire net_2541;
wire net_391;
wire net_1002;
wire net_533;
wire net_2297;
wire net_3325;
wire net_1695;
wire net_911;
wire net_1617;
wire x1214;
wire net_3188;
wire net_37;
wire net_2048;
wire net_582;
wire net_2341;
wire net_1993;
wire net_3010;
wire net_661;
wire net_881;
wire net_3360;
wire net_2805;
wire net_2903;
wire net_2516;
wire net_1397;
wire net_568;
wire net_2807;
wire net_47;
wire net_1141;
wire net_1227;
wire net_3243;
wire net_1008;
wire net_1543;
wire net_1295;
wire net_2104;
wire net_1954;
wire net_1443;
wire net_1288;
wire net_3069;
wire net_3170;
wire net_2071;
wire net_2840;
wire net_1923;
wire net_1275;
wire net_210;
wire net_2766;
wire net_2155;
wire net_168;
wire net_2417;
wire net_2300;
wire net_2041;
wire net_916;
wire net_3395;
wire net_3199;
wire net_741;
wire net_940;
wire net_385;
wire net_2609;
wire net_851;
wire net_269;
wire net_3193;
wire net_3131;
wire net_469;
wire net_2426;
wire net_3179;
wire net_1978;
wire net_1945;
wire net_3167;
wire net_1170;
wire x597;
wire net_2423;
wire net_1833;
wire net_3310;
wire net_1043;
wire net_671;
wire net_2280;
wire net_2831;
wire net_3029;
wire net_2850;
wire net_2366;
wire net_778;
wire net_2380;
wire net_3393;
wire net_770;
wire net_2930;
wire net_1455;
wire net_1005;
wire x1427;
wire net_1059;
wire net_1630;
wire net_895;
wire net_1454;
wire net_2956;
wire x1186;
wire net_307;
wire net_1796;
wire net_1082;
wire net_3342;
wire net_1412;
wire net_1550;
wire net_2310;
wire net_1507;
wire net_3296;
wire net_257;
wire net_233;
wire net_1255;
wire net_474;
wire net_2656;
wire net_958;
wire x1980;
wire net_1250;
wire net_1481;
wire net_1268;
wire net_995;
wire net_3212;
wire x808;
wire net_3040;
wire net_1115;
wire net_207;
wire net_944;
wire net_1734;
wire net_1764;
wire net_700;
wire net_961;
wire net_1246;
wire net_3004;
wire net_2106;
wire net_3335;
wire x49;
wire net_1689;
wire net_1774;
wire net_3050;
wire net_1728;
wire net_1673;
wire net_63;
wire net_3327;
wire net_3060;
wire net_2667;
wire net_274;
wire net_2568;
wire x935;
wire net_1075;
wire net_321;
wire net_425;
wire net_287;
wire net_189;
wire net_2387;
wire net_1586;
wire net_930;
wire net_833;
wire net_2995;
wire net_2205;
wire net_99;
wire net_2945;
wire net_480;
wire x663;
wire net_2267;
wire net_216;
wire net_934;
wire net_2897;
wire net_433;
wire net_3103;
wire net_2881;
wire net_836;
wire net_544;
wire net_717;
wire net_2161;
wire x956;
wire net_368;
wire net_224;
wire net_1399;
wire net_52;
wire net_1898;
wire net_1824;
wire net_608;
wire net_1212;
wire net_3350;
wire net_370;
wire net_3402;
wire net_2223;
wire net_2000;
wire net_2673;
wire x990;
wire net_2984;
wire net_1120;
wire net_1020;
wire net_2848;
wire net_3166;
wire net_3282;
wire net_3304;
wire net_3122;
wire net_1169;
wire net_973;
wire net_1139;
wire net_1245;
wire net_2549;
wire net_2206;
wire net_1781;
wire net_860;
wire net_1392;
wire net_870;
wire net_1574;
wire net_3049;
wire net_2046;
wire net_2094;
wire net_2543;
wire net_637;
wire net_311;
wire net_2878;
wire net_760;
wire net_2871;
wire net_2514;
wire net_2479;
wire net_2083;
wire net_2390;
wire net_873;
wire net_2488;
wire net_1811;
wire net_154;
wire net_3267;
wire net_2321;
wire net_2686;
wire net_2013;
wire net_2588;
wire net_1509;
wire net_817;
wire net_1870;
wire net_529;
wire net_3414;
wire net_704;
wire net_2520;
wire net_1478;
wire net_2179;
wire net_1696;
wire net_587;
wire net_1262;
wire net_97;
wire net_2028;
wire net_2553;
wire net_2063;
wire net_192;
wire net_1889;
wire net_1739;
wire net_1356;
wire net_2912;
wire x1014;
wire net_2920;
wire net_2197;
wire net_1591;
wire x1073;
wire x870;
wire net_2981;
wire x166;
wire net_1747;
wire net_2012;
wire net_1164;
wire net_650;
wire net_735;
wire net_2905;
wire net_1907;
wire net_121;
wire net_1711;
wire net_200;
wire net_597;
wire net_2084;
wire net_743;
wire net_2583;
wire net_1922;
wire net_195;
wire net_1081;
wire net_1853;
wire net_2037;
wire net_2170;
wire x1710;
wire net_2664;
wire net_1237;
wire net_1420;
wire net_2706;
wire net_849;
wire net_2678;
wire net_603;
wire x444;
wire net_2451;
wire net_2602;
wire net_401;
wire net_642;
wire net_2699;
wire net_1522;
wire net_1158;
wire net_3144;
wire net_2926;
wire net_2714;
wire net_699;
wire net_242;
wire net_2183;
wire net_2557;
wire net_359;
wire net_440;
wire net_2526;
wire x152;
wire net_470;
wire net_758;
wire net_2702;
wire net_2819;
wire net_1644;
wire net_430;
wire net_2864;
wire net_2834;
wire net_2800;
wire net_882;
wire net_718;
wire net_1998;
wire x64;
wire net_1827;
wire net_3225;
wire net_1190;
wire net_83;
wire net_2795;
wire x144;
wire net_1311;
wire net_3129;
wire net_2283;
wire net_1207;
wire net_3255;
wire net_1918;
wire net_56;
wire x850;
wire net_2121;
wire net_1063;
wire net_2191;
wire net_968;
wire x1456;
wire net_336;
wire net_3236;
wire net_3201;
wire net_2252;
wire net_555;
wire net_1578;
wire net_2534;
wire net_1613;
wire net_2917;
wire net_3221;
wire net_790;
wire net_2126;
wire net_1504;
wire net_697;
wire net_2003;
wire net_475;
wire net_1577;
wire net_1417;
wire net_1054;
wire net_3411;
wire net_605;
wire x0;
wire net_2309;
wire net_2386;
wire net_2727;
wire net_2166;
wire net_502;
wire net_2470;
wire net_2465;
wire net_1564;
wire net_2257;
wire net_1568;
wire net_3418;
wire net_2304;
wire x629;
wire net_924;
wire net_1526;
wire net_898;
wire net_2968;
wire net_1884;
wire net_1333;
wire net_2643;
wire net_2348;
wire net_1593;
wire net_489;
wire net_2646;
wire net_3082;
wire net_714;
wire net_2999;
wire net_1309;
wire net_3380;
wire net_683;
wire net_1771;
wire net_148;
wire net_1376;
wire net_2628;
wire net_2748;
wire net_1517;
wire net_1980;
wire net_1360;
wire net_251;
wire net_2054;
wire net_3364;
wire net_1302;
wire net_2076;
wire net_244;
wire net_2218;
wire net_664;
wire net_128;
wire net_840;
wire net_2395;
wire net_1690;
wire net_1364;
wire net_1078;
wire net_549;
wire net_827;
wire net_1989;
wire net_2997;
wire net_2855;
wire net_2793;
wire net_2093;
wire net_1795;
wire net_411;
wire net_2137;
wire net_1836;
wire x245;
wire net_2337;
wire net_2403;
wire net_1539;
wire net_1369;
wire x136;
wire net_1862;
wire net_2317;
wire x2116;
wire x730;
wire net_3035;
wire net_2355;
wire net_1013;
wire net_1530;
wire net_3075;
wire net_3262;
wire net_2952;
wire net_1548;
wire net_842;
wire net_92;
wire net_112;
wire net_394;
wire net_810;
wire net_2336;
wire net_1705;
wire net_2536;
wire net_1189;
wire net_139;
wire net_2035;
wire net_2373;
wire net_409;
wire net_2949;
wire net_2826;
wire net_1469;
wire net_2398;
wire net_492;
wire net_88;
wire net_2141;
wire net_1708;
wire net_2639;
wire net_2436;
wire net_3315;
wire x701;
wire net_81;
wire net_2455;
wire net_1609;
wire net_402;
wire net_1327;
wire net_110;
wire net_3419;
wire net_2976;
wire net_722;
wire net_33;
wire net_1403;
wire net_3248;
wire net_988;
wire net_1254;
wire net_2248;
wire net_2274;
wire net_2270;
wire net_1667;
wire net_621;
wire net_435;
wire net_1606;
wire net_1386;
wire x397;
wire net_1830;
wire net_2359;
wire net_132;
wire net_105;
wire net_2838;
wire net_3054;
wire net_1649;
wire net_1837;
wire net_1841;
wire net_1249;
wire net_2427;
wire net_3378;
wire net_1071;
wire net_2186;
wire net_3163;
wire net_2868;
wire net_2029;
wire net_1430;
wire net_569;
wire net_2478;
wire net_2563;
wire net_2946;
wire net_327;
wire net_2587;
wire net_3408;
wire net_1284;
wire net_1701;
wire net_630;
wire net_2959;
wire net_999;
wire net_76;
wire net_2202;
wire net_1888;
wire net_2490;
wire x1681;
wire net_353;
wire net_822;
wire net_1633;
wire net_1791;
wire net_1471;
wire net_1792;
wire net_2496;
wire net_3109;
wire net_2066;
wire net_1974;
wire net_1480;
wire net_319;
wire net_2670;
wire net_1743;
wire net_1598;
wire net_3124;
wire net_3046;
wire net_2597;
wire net_1903;
wire net_164;
wire net_2407;
wire x692;
wire net_377;
wire net_731;
wire net_1146;
wire net_87;
wire net_1544;
wire net_288;
wire net_912;
wire net_2649;
wire net_3096;
wire net_1629;
wire net_1459;
wire net_3277;
wire net_805;
wire x1844;
wire net_1733;
wire net_2923;
wire net_2151;
wire net_2078;
wire net_540;
wire net_512;
wire net_779;
wire net_2688;
wire net_2642;
wire net_1928;
wire net_1174;
wire net_1622;
wire net_891;
wire x98;
wire net_1328;
wire net_1109;
wire net_234;
wire net_2859;
wire net_38;
wire net_3065;
wire net_2884;
wire net_3102;
wire net_2762;
wire net_3205;
wire net_1102;
wire net_1094;
wire net_2749;
wire net_1724;
wire net_855;
wire net_674;
wire net_3371;
wire net_618;
wire net_2244;
wire net_2692;
wire x83;
wire net_303;
wire net_2089;
wire net_2475;
wire net_1875;
wire net_491;
wire net_965;
wire x1582;
wire net_1299;
wire x1110;
wire net_3420;
wire net_2937;
wire net_948;
wire net_783;
wire net_1487;
wire net_1195;
wire net_2916;
wire net_754;
wire net_2759;
wire x355;
wire net_421;
wire net_2502;
wire net_1396;
wire net_2605;
wire net_1104;
wire net_921;
wire net_550;
wire net_764;
wire net_2593;
wire net_876;
wire net_2737;
wire net_2162;
wire net_2439;
wire net_3308;
wire net_172;
wire net_2481;
wire net_2835;
wire net_2192;
wire net_1533;
wire net_1117;
wire net_1458;
wire net_1240;
wire net_461;
wire net_3000;
wire net_2564;
wire net_905;
wire net_2617;
wire net_1060;
wire net_2821;
wire net_1512;
wire net_1658;
wire net_142;
wire net_654;
wire net_858;
wire net_330;
wire net_2235;
wire net_2229;
wire net_1330;
wire net_158;
wire net_3200;
wire net_1715;
wire net_3007;
wire net_2080;
wire net_3015;
wire net_1785;
wire net_2711;
wire net_2097;
wire net_3174;
wire x1170;
wire net_2876;
wire net_2504;
wire net_570;
wire net_444;
wire net_525;
wire net_844;
wire net_2175;
wire net_1496;
wire net_1216;
wire net_1210;
wire net_1067;
wire net_325;
wire net_2815;
wire net_1820;
wire x1769;
wire net_1427;
wire net_1271;
wire net_1086;
wire net_2116;
wire net_1758;
wire x1863;
wire net_985;
wire net_1782;
wire net_1769;
wire net_1197;
wire net_1967;
wire net_1278;
wire net_273;
wire net_424;
wire net_1567;
wire net_3182;
wire net_576;
wire net_1654;
wire net_1521;
wire x78;
wire net_1729;
wire net_3353;
wire net_2098;
wire net_1677;
wire net_465;
wire net_3355;
wire net_177;
wire net_3005;
wire net_1883;
wire net_2991;
wire net_2783;
wire net_476;
wire net_564;
wire net_2803;
wire net_2050;
wire net_382;
wire net_3301;
wire net_3058;
wire net_725;
wire net_2811;
wire net_3086;
wire net_1315;
wire net_583;
wire net_2058;
wire net_813;
wire net_3045;
wire net_1178;
wire net_953;
wire net_2612;
wire net_1027;
wire net_894;
wire net_1074;
wire net_2018;
wire net_1058;
wire x44;
wire net_1423;
wire net_2042;
wire net_340;
wire net_2902;
wire net_1871;
wire net_1408;
wire net_2510;
wire net_265;
wire net_517;
wire net_2634;
wire net_434;
wire net_628;
wire net_2489;
wire net_1465;
wire net_220;
wire net_1797;
wire net_293;
wire x1636;
wire net_3023;
wire net_1202;
wire net_1938;
wire net_69;
wire net_543;
wire x201;
wire net_1155;
wire net_3160;
wire net_925;
wire net_2125;
wire net_625;
wire net_339;
wire net_2279;
wire net_1823;
wire net_2695;
wire net_864;
wire x331;
wire net_1289;
wire net_3138;
wire net_2623;
wire net_261;
wire net_191;
wire net_2909;
wire net_2710;
wire net_558;
wire net_2069;
wire x1318;
wire net_2660;
wire net_2362;
wire net_2298;
wire net_660;
wire net_1618;
wire net_102;
wire net_2313;
wire net_59;
wire net_2497;
wire net_1955;
wire net_2723;
wire net_2552;
wire net_1908;
wire x295;
wire net_3229;
wire net_1001;
wire net_3217;
wire net_1694;
wire net_781;
wire net_1291;
wire net_230;
wire net_1865;
wire net_910;
wire x1047;
wire net_3383;
wire net_678;
wire net_3012;
wire net_3349;
wire net_2412;
wire net_185;
wire net_1222;
wire net_3404;
wire net_928;
wire net_1984;
wire net_2578;
wire net_208;
wire net_1994;
wire net_1375;
wire net_1015;
wire net_315;
wire net_2980;
wire net_2744;
wire net_2377;
wire net_1944;
wire net_1433;
wire net_415;
wire net_1351;
wire net_116;
wire net_1775;
wire net_3251;
wire net_2786;
wire net_347;
wire net_1535;
wire net_297;
wire net_91;
wire net_346;
wire net_2400;
wire net_3358;
wire net_1776;
wire net_2287;
wire net_2145;
wire net_448;
wire net_3368;
wire net_2034;
wire net_1335;
wire net_2574;
wire net_886;
wire net_229;
wire net_3311;
wire net_3189;
wire net_1808;
wire net_3256;
wire net_2988;
wire net_2146;
wire net_687;
wire net_3266;
wire net_2212;
wire net_405;
wire net_2132;
wire net_2292;
wire net_1111;
wire x1719;
wire net_2651;
wire net_1880;
wire net_184;
wire net_3322;
wire net_3155;
wire net_2533;
wire net_610;
wire net_1844;
wire net_1470;
wire net_1913;
wire net_389;
wire x1877;
wire net_831;
wire net_902;
wire net_1867;
wire net_451;
wire net_2344;
wire net_1323;
wire net_2650;
wire net_1949;
wire net_1506;
wire x2167;
wire x543;
wire net_1234;
wire net_750;
wire net_1583;
wire net_736;
wire net_1804;
wire net_1760;
wire net_539;
wire net_2331;
wire net_692;
wire net_1184;
wire net_1563;
wire net_2778;
wire net_2756;
wire net_3361;
wire net_1365;
wire net_1135;
wire net_1346;
wire net_43;
wire net_3403;
wire net_1960;
wire net_1085;
wire x229;
wire net_1942;
wire net_592;
wire net_3093;
wire net_1801;
wire net_3247;
wire net_1400;
wire net_647;
wire net_885;
wire net_1267;
wire net_773;
wire net_2464;
wire net_2266;
wire net_281;
wire x1993;
wire net_828;
wire net_869;
wire net_1603;
wire x57;
wire net_669;
wire net_2732;
wire net_937;
wire net_2441;
wire x574;
wire x484;
wire net_2349;
wire net_496;
wire net_761;
wire net_1554;
wire net_479;
wire net_1096;
wire net_1294;
wire net_795;
wire net_982;
wire net_2459;
wire net_2030;
wire net_1587;
wire net_1354;
wire net_1580;
wire net_2904;
wire net_796;
wire net_1308;
wire net_1406;
wire net_2249;
wire net_54;
wire net_526;
wire net_2718;
wire net_834;
wire net_694;
wire net_648;
wire net_1389;
wire net_2747;
wire net_739;
wire net_1434;
wire net_974;
wire net_1570;
wire net_3250;
wire x1361;
wire net_774;
wire net_2548;
wire net_2075;
wire net_826;
wire net_923;
wire net_1738;
wire net_548;
wire net_3359;
wire net_2402;
wire net_1707;
wire net_2190;
wire net_1881;
wire net_501;
wire x621;
wire net_111;
wire net_2624;
wire net_225;
wire net_636;
wire net_124;
wire net_252;
wire net_343;
wire net_3323;
wire net_3128;
wire net_2399;
wire net_511;
wire net_901;
wire net_1961;
wire net_447;
wire net_2611;
wire net_871;
wire net_1260;
wire net_3425;
wire net_410;
wire net_2654;
wire net_390;
wire net_1492;
wire net_2487;
wire net_35;
wire net_2911;
wire net_1154;
wire net_1185;
wire net_1819;
wire x121;
wire net_2537;
wire net_239;
wire net_310;
wire net_2975;
wire net_2437;
wire net_2779;
wire x1466;
wire net_80;
wire net_1912;
wire net_2951;
wire net_2603;
wire net_1132;
wire net_1490;
wire net_2442;
wire net_2293;
wire net_682;
wire net_280;
wire net_989;
wire net_1963;
wire x1750;
wire net_1538;
wire net_3026;
wire net_495;
wire net_34;
wire net_108;
wire net_458;
wire x857;
wire net_685;
wire net_1802;
wire net_2356;
wire net_2140;
wire net_3288;
wire net_971;
wire x253;
wire net_2273;
wire net_2049;
wire net_617;
wire net_2517;
wire net_2316;
wire net_2184;
wire net_554;
wire net_1007;
wire net_1579;
wire net_1292;
wire net_2755;
wire net_1999;
wire net_1014;
wire net_2703;
wire net_1678;
wire net_2796;
wire net_46;
wire net_1444;
wire net_2679;
wire net_3366;
wire net_584;
wire net_1441;
wire net_3410;
wire net_2111;
wire net_1946;
wire net_2733;
wire net_969;
wire net_1525;
wire net_2411;
wire x1063;
wire net_165;
wire net_538;
wire net_1605;
wire net_1937;
wire net_821;
wire net_2535;
wire net_3191;
wire net_366;
wire net_1956;
wire net_1854;
wire net_1917;
wire net_1614;
wire net_1755;
wire net_747;
wire net_1359;
wire net_2305;
wire net_1653;
wire net_2335;
wire net_2460;
wire net_2983;
wire net_3209;
wire net_384;
wire x1915;
wire net_2258;
wire net_198;
wire net_1647;
wire net_2618;
wire net_3365;
wire net_209;
wire net_1282;
wire x1368;
wire net_294;
wire net_2599;
wire net_2665;
wire net_2367;
wire net_2892;
wire net_2707;
wire net_1114;
wire net_2810;
wire net_2429;
wire net_3204;
wire net_1265;
wire net_3388;
wire net_1053;
wire net_1004;
wire net_485;
wire net_848;
wire net_1748;
wire net_3078;
wire net_3218;
wire net_1080;
wire net_1619;
wire net_3232;
wire net_2124;
wire net_2964;
wire net_1890;
wire net_1161;
wire x36;
wire net_3334;
wire net_3224;
wire net_82;
wire net_64;
wire net_3228;
wire net_2343;
wire net_2232;
wire net_1719;
wire net_2282;
wire net_726;
wire net_2430;
wire net_2357;
wire net_1028;
wire net_1529;
wire net_600;
wire net_3237;
wire net_1395;
wire net_1546;
wire net_701;
wire net_125;
wire net_397;
wire x159;
wire net_808;
wire net_1589;
wire net_1046;
wire net_2440;
wire net_1685;
wire net_1704;
wire net_606;
wire net_623;
wire net_2396;
wire net_663;
wire net_1213;
wire net_1384;
wire net_2738;
wire net_1891;
wire net_1379;
wire net_2265;
wire net_320;
wire net_1322;
wire net_579;
wire net_2445;
wire net_2644;
wire net_2944;
wire net_769;
wire net_3396;
wire net_1301;
wire net_1780;
wire net_2062;
wire net_986;
wire net_1242;
wire net_2856;
wire net_286;
wire x1800;
wire net_787;
wire net_1241;
wire x459;
wire net_2894;
wire net_1025;
wire net_1988;
wire net_935;
wire net_3001;
wire x523;
wire net_3116;
wire net_1511;
wire net_645;
wire net_1518;
wire net_3121;
wire net_426;
wire net_1089;
wire net_1194;
wire net_1437;
wire net_1634;
wire net_414;
wire net_609;
wire x1662;
wire net_1048;
wire net_1664;
wire net_3048;
wire net_799;
wire net_3083;
wire net_705;
wire net_2139;
wire x585;
wire net_1608;
wire net_506;
wire net_2948;
wire net_1816;
wire net_2014;
wire net_1910;
wire net_1221;
wire net_1036;
wire net_1951;
wire x554;
wire net_331;
wire net_3034;
wire net_1196;
wire net_816;
wire net_3264;
wire net_2493;
wire net_919;
wire net_2558;
wire net_2092;
wire net_2454;
wire net_2220;
wire net_2040;
wire net_2823;
wire net_290;
wire net_1217;
wire net_1508;
wire net_3379;
wire net_3313;
wire net_3136;
wire net_2933;
wire net_931;
wire net_3381;
wire net_2209;
wire x1645;
wire net_1372;
wire net_1757;
wire net_2242;
wire x2143;
wire x675;
wire net_759;
wire net_1575;
wire net_3279;
wire x1593;
wire net_3152;
wire net_2682;
wire net_657;
wire net_1727;
wire net_140;
wire net_247;
wire net_740;
wire net_329;
wire net_1722;
wire net_2329;
wire net_2150;
wire net_2008;
wire net_1259;
wire net_2065;
wire x185;
wire net_1924;
wire net_2839;
wire net_2143;
wire net_1825;
wire net_3183;
wire net_2927;
wire net_2196;
wire net_3413;
wire net_3168;
wire net_70;
wire net_2808;
wire net_194;
wire net_2178;
wire net_730;
wire net_962;
wire net_1341;
wire net_478;
wire net_1934;
wire net_3242;
wire net_1128;
wire net_1835;
wire net_3073;
wire net_2713;
wire net_2105;
wire net_596;
wire net_1127;
wire net_1848;
wire net_1261;
wire net_333;
wire net_804;
wire net_639;
wire net_1119;
wire net_2120;
wire net_1975;
wire net_1314;
wire net_957;
wire net_1287;
wire net_1238;
wire net_2726;
wire net_531;
wire net_2569;
wire net_77;
wire net_499;
wire net_565;
wire net_3345;
wire net_2752;
wire x2062;
wire net_2832;
wire net_49;
wire net_1033;
wire net_1340;
wire net_3028;
wire net_2149;
wire net_3123;
wire net_2955;
wire net_2554;
wire net_71;
wire net_3328;
wire net_1692;
wire net_771;
wire net_2655;
wire net_2528;
wire x1868;
wire net_1765;
wire net_2844;
wire net_2301;
wire net_3107;
wire net_2978;
wire net_2107;
wire x1933;
wire net_1686;
wire net_180;
wire net_1361;
wire net_367;
wire net_3303;
wire net_51;
wire net_2774;
wire net_2420;
wire net_2450;
wire net_2860;
wire net_432;
wire net_1979;
wire net_1062;
wire net_1842;
wire net_1208;
wire net_3290;
wire net_3293;
wire net_204;
wire net_1142;
wire net_1460;
wire net_1475;
wire net_1451;
wire net_232;
wire net_3159;
wire net_67;
wire net_2240;
wire net_1180;
wire net_2416;
wire net_1627;
wire net_2002;
wire net_1069;
wire net_2022;
wire net_2167;
wire net_2880;
wire net_203;
wire net_1411;
wire net_2385;
wire net_2173;
wire net_2996;
wire net_505;
wire net_2889;
wire net_1602;
wire net_137;
wire net_1416;
wire net_992;
wire net_237;
wire net_613;
wire net_3154;
wire net_2433;
wire net_782;
wire net_2144;
wire net_2501;
wire net_532;
wire net_2236;
wire net_93;
wire net_1601;
wire net_2729;
wire net_1916;
wire net_1095;
wire net_578;
wire net_3314;
wire net_2971;
wire net_2468;
wire x216;
wire net_302;
wire net_1131;
wire net_889;
wire net_1116;
wire net_348;
wire net_1558;
wire net_753;
wire net_2743;
wire net_2836;
wire net_1505;
wire net_626;
wire net_1805;
wire net_2159;
wire net_388;
wire x1262;
wire net_100;
wire net_1809;
wire net_1861;
wire net_2195;
wire net_536;
wire net_686;
wire net_455;
wire net_1615;
wire net_1332;
wire net_3421;
wire net_2814;
wire net_221;
wire net_1594;
wire net_115;
wire x114;
wire net_1691;
wire net_3339;
wire net_3276;
wire net_689;
wire net_1110;
wire net_393;
wire net_751;
wire net_442;
wire net_2112;
wire net_542;
wire net_595;
wire net_2363;
wire net_408;
wire net_1832;
wire net_1320;
wire net_1026;
wire net_1828;
wire net_3246;
wire net_2215;
wire net_1466;
wire net_1845;
wire net_2573;
wire net_3087;
wire net_2376;
wire net_1520;
wire net_157;
wire x302;
wire net_1710;
wire net_1821;
wire net_42;
wire net_1228;
wire net_1205;
wire net_3390;
wire net_1401;
wire net_2372;
wire net_1588;
wire net_66;
wire net_466;
wire net_868;
wire net_1179;
wire net_1495;
wire net_2722;
wire net_2992;
wire net_1426;
wire net_3039;
wire net_3233;
wire net_2217;
wire net_3147;
wire net_938;
wire net_1407;
wire net_443;
wire net_1610;
wire net_1761;
wire net_270;
wire net_522;
wire net_922;
wire net_3263;
wire net_183;
wire net_2638;
wire net_668;
wire net_1440;
wire net_3079;
wire net_1057;
wire net_2915;
wire net_1584;
wire net_1990;
wire net_1011;
wire net_2330;
wire net_1355;
wire net_2264;
wire net_800;
wire net_644;
wire net_977;
wire net_643;
wire net_3397;
wire net_1070;
wire net_852;
wire net_2987;
wire net_1225;
wire net_622;
wire net_812;
wire net_2253;
wire net_2580;
wire x1958;
wire net_1699;
wire net_1042;
wire net_1385;
wire net_1643;
wire net_2857;
wire net_1107;
wire net_1919;
wire net_1534;
wire net_2767;
wire x899;
wire net_1000;
wire net_1338;
wire net_2045;
wire net_2521;
wire net_2053;
wire net_1995;
wire net_2545;
wire net_3384;
wire net_1016;
wire net_2180;
wire net_1203;
wire net_2869;
wire net_3332;
wire net_825;
wire net_1892;
wire net_1798;
wire net_3220;
wire net_2119;
wire net_309;
wire net_659;
wire x883;
wire net_29;
wire net_1366;
wire net_837;
wire net_2615;
wire x1554;
wire net_899;
wire net_1744;
wire net_516;
wire net_1010;
wire net_2870;
wire net_31;
wire net_1693;
wire net_3176;
wire net_927;
wire net_2007;
wire net_956;
wire net_1151;
wire net_2908;
wire net_2068;
wire net_713;
wire net_693;
wire net_1519;
wire net_2596;
wire x2080;
wire net_729;
wire net_2970;
wire net_3213;
wire net_2818;
wire net_863;
wire x638;
wire net_2675;
wire net_438;
wire net_2794;
wire net_3164;
wire net_2584;
wire net_580;
wire net_314;
wire net_1752;
wire net_2250;
wire net_2136;
wire net_904;
wire net_2527;
wire net_2339;
wire net_3013;
wire net_341;
wire net_3110;
wire net_952;
wire net_2967;
wire net_2091;
wire net_2406;
wire net_58;
wire net_1879;
wire net_3185;
wire net_970;
wire net_488;
wire net_3300;
wire net_807;
wire net_3405;
wire net_3270;
wire net_86;
wire x1333;
wire net_2319;
wire net_2245;
wire net_3044;
wire net_1532;
wire net_2474;
wire net_1160;
wire net_945;
wire net_2530;
wire net_159;
wire net_2101;
wire net_3268;
wire net_2163;
wire net_383;
wire net_3417;
wire net_3307;
wire x815;
wire net_217;
wire net_553;
wire net_3140;
wire net_1093;
wire net_2592;
wire x128;
wire net_2875;
wire net_427;
wire net_763;
wire net_2785;
wire net_135;
wire net_915;
wire net_3259;
wire net_2226;
wire net_1121;
wire net_473;
wire net_1740;
wire net_324;
wire net_710;
wire net_2777;
wire net_1049;
wire net_454;
wire net_418;
wire net_462;
wire net_872;
wire net_1784;
wire net_3097;
wire net_1296;
wire net_161;
wire net_709;
wire net_2484;
wire net_2863;
wire net_3066;
wire net_1066;
wire net_1165;
wire net_677;
wire net_3018;
wire net_2606;
wire net_173;
wire net_1472;
wire net_1486;
wire net_2939;
wire net_78;
wire net_2424;
wire net_1113;
wire net_2591;
wire net_2320;
wire net_1968;
wire net_1839;
wire net_1665;
wire net_1344;
wire net_3006;
wire net_376;
wire net_1084;
wire net_1283;
wire net_354;
wire net_1500;
wire net_2133;
wire net_1681;
wire x535;
wire net_2507;
wire net_1136;
wire net_2515;
wire net_1812;
wire net_3173;
wire net_3008;
wire net_2685;
wire net_2763;
wire net_2898;
wire net_2658;
wire net_573;
wire net_2174;
wire net_1391;
wire net_3356;
wire net_2224;
wire net_784;
wire net_3203;
wire net_422;
wire net_1772;
wire net_1345;
wire net_1450;
wire net_561;
wire net_45;
wire net_2659;
wire net_2589;
wire net_2498;
wire net_381;
wire net_591;
wire net_1700;
wire net_746;
wire net_2326;
wire net_1592;
wire net_2085;
wire net_2290;
wire net_1274;
wire net_2458;
wire net_1682;
wire net_2851;
wire net_178;
wire net_1857;
wire net_2843;
wire net_2635;
wire net_1637;
wire net_3374;
wire x562;
wire net_3238;
wire net_1318;
wire net_2698;
wire net_941;
wire net_809;
wire net_629;
wire net_1663;
wire net_55;
wire net_1557;
wire net_635;
wire net_266;
wire net_1235;
wire net_2691;
wire net_1037;
wire net_1514;
wire net_2019;
wire net_3092;
wire x439;
wire net_2311;
wire net_2070;
wire net_350;
wire net_3019;
wire x1031;
wire net_1599;
wire net_306;
wire net_2351;
wire net_3132;
wire net_3161;
wire net_3117;
wire net_1290;
wire net_500;
wire net_1350;
wire net_3053;
wire net_1906;
wire net_3198;
wire net_2610;
wire x1611;
wire net_1626;
wire net_1648;
wire net_2822;
wire net_1258;
wire net_2982;
wire net_1623;
wire net_631;
wire x467;
wire net_3297;
wire net_2023;
wire net_3369;
wire net_123;
wire net_1329;
wire x347;
wire net_1101;
wire net_994;
wire net_262;
wire net_362;
wire net_527;
wire net_1668;
wire net_3424;
wire net_3127;
wire net_318;
wire net_1052;
wire net_1971;
wire net_3139;
wire net_2409;
wire net_3192;
wire net_1900;
wire net_1793;
wire net_1779;
wire net_3104;
wire net_2647;
wire net_670;
wire net_2189;
wire net_2278;
wire net_2057;
wire net_3340;
wire net_3072;
wire net_103;
wire net_226;
wire net_1124;
wire net_2687;
wire net_1849;
wire net_1021;
wire net_228;
wire net_1737;
wire net_2640;
wire net_143;
wire net_966;
wire net_1859;
wire net_3372;
wire net_190;
wire net_2887;
wire net_1447;
wire net_1920;
wire net_145;
wire net_2201;
wire net_1929;
wire net_1108;
wire net_2827;
wire net_2025;
wire net_2010;
wire net_1983;
wire x413;
wire net_2936;
wire net_3030;
wire net_2061;
wire net_1145;
wire net_2804;
wire net_1878;
wire net_2261;
wire net_188;
wire net_1553;
wire net_3061;
wire net_1895;
wire net_3319;
wire net_509;
wire net_755;
wire x389;
wire net_1723;
wire net_2491;
wire net_211;
wire net_2900;
wire net_133;
wire net_2958;
wire net_3208;
wire net_1077;
wire net_2924;
wire net_2704;
wire net_3151;
wire net_2410;
wire net_2306;
wire net_1851;
wire x451;
wire net_3272;
wire net_2873;
wire net_557;
wire net_3108;
wire net_119;
wire net_3043;
wire net_2254;
wire x761;
wire net_2861;
wire net_2185;
wire net_1652;
wire net_2669;
wire net_2233;
wire net_1321;
wire net_1429;
wire net_2941;
wire net_2033;
wire x378;
wire net_3348;
wire net_1991;
wire net_477;
wire net_1611;
wire net_2123;
wire net_1173;
wire net_1209;
wire net_1431;
wire net_1754;
wire net_2725;
wire net_1099;
wire net_2328;
wire net_2943;
wire x1517;
wire net_1714;
wire net_2532;
wire net_727;
wire net_847;
wire net_90;
wire net_2315;
wire net_283;
wire net_2231;
wire net_85;
wire x1490;
wire net_3190;
wire net_1864;
wire net_404;
wire net_240;
wire net_1200;
wire net_2518;
wire net_2666;
wire net_295;
wire net_1239;
wire net_1463;
wire net_344;
wire net_2269;
wire net_884;
wire net_1646;
wire net_712;
wire net_2281;
wire net_1422;
wire net_2776;
wire net_2259;
wire net_2056;
wire net_3389;
wire x1808;
wire net_1562;
wire net_2522;
wire net_472;
wire net_1106;
wire net_65;
wire net_1510;
wire net_1628;
wire net_1394;
wire net_2963;
wire net_3077;
wire net_2972;
wire net_2739;
wire x421;
wire net_484;
wire net_896;
wire net_1281;
wire net_2512;
wire net_2110;
wire net_3223;
wire net_2463;
wire net_2919;
wire net_136;
wire net_1936;
wire net_1524;
wire net_2893;
wire net_2241;
wire net_3227;
wire net_2358;
wire net_1528;
wire net_126;
wire net_2708;
wire net_278;
wire net_1749;
wire net_3367;
wire net_3057;
wire x273;
wire net_1547;
wire net_2211;
wire net_571;
wire net_601;
wire net_1162;
wire net_1362;
wire net_1896;
wire net_2443;
wire net_2472;
wire net_1307;
wire net_2346;
wire net_2790;
wire net_2742;
wire net_1982;
wire net_1732;
wire net_2511;
wire net_1877;
wire net_829;
wire net_2626;
wire x237;
wire net_720;
wire net_2294;
wire net_2115;
wire net_2299;
wire net_2393;
wire net_2199;
wire net_3376;
wire net_900;
wire net_3320;
wire net_1405;
wire net_2625;
wire net_684;
wire net_3253;
wire net_2648;
wire net_1882;
wire net_510;
wire net_1353;
wire net_413;
wire net_1595;
wire net_2001;
wire net_1491;
wire net_716;
wire net_114;
wire net_1269;
wire net_2653;
wire net_2419;
wire net_1300;
wire x515;
wire net_2974;
wire net_2960;
wire net_1034;
wire net_36;
wire net_1252;
wire net_2696;
wire net_2734;
wire net_253;
wire net_276;
wire net_2782;
wire net_494;
wire net_1449;
wire x506;
wire net_547;
wire x1835;
wire net_1098;
wire net_666;
wire net_3146;
wire net_507;
wire net_1959;
wire net_1902;
wire net_616;
wire net_238;
wire net_1220;
wire net_28;
wire net_3074;
wire net_1847;
wire net_2438;
wire net_2600;
wire net_1911;
wire net_3022;
wire net_2717;
wire net_793;
wire net_649;
wire net_460;
wire net_1657;
wire net_3084;
wire x106;
wire net_1374;
wire net_2353;
wire net_1962;
wire net_457;
wire net_291;
wire net_2246;
wire net_2272;
wire net_1964;
wire net_772;
wire net_2494;
wire net_857;
wire net_867;
wire net_2334;
wire net_1367;
wire net_396;
wire net_1133;
wire net_3287;
wire net_166;
wire net_107;
wire net_1277;
wire net_2866;
wire net_1976;
wire net_2661;
wire net_3169;
wire net_530;
wire net_1541;
wire net_3025;
wire x1244;
wire net_1371;
wire net_3352;
wire net_2758;
wire net_594;
wire net_271;
wire net_3329;
wire net_117;
wire net_74;
wire net_673;
wire net_1826;
wire net_2064;
wire net_205;
wire net_1286;
wire net_2797;
wire net_2852;
wire net_1721;
wire net_1925;
wire x748;
wire net_2142;
wire net_1445;
wire net_2074;
wire net_1909;
wire net_920;
wire net_1952;
wire net_334;
wire net_2577;
wire net_1410;
wire net_2954;
wire net_1461;
wire net_3062;
wire net_3009;
wire net_2453;
wire net_1073;
wire net_365;
wire net_3274;
wire net_1947;
wire net_3177;
wire net_820;
wire net_3344;
wire net_2953;
wire net_380;
wire net_2847;
wire net_141;
wire net_467;
wire net_879;
wire net_1810;
wire net_1118;
wire net_2910;
wire net_1556;
wire net_2415;
wire net_372;
wire net_2990;
wire net_2081;
wire net_437;
wire x1286;
wire net_1270;
wire net_2286;
wire net_566;
wire net_1552;
wire net_803;
wire net_3165;
wire x434;
wire net_3197;
wire net_2788;
wire net_624;
wire net_1348;
wire net_2148;
wire x20;
wire net_1476;
wire net_3215;
wire net_2108;
wire net_1933;
wire net_298;
wire net_1293;
wire net_2529;
wire net_688;
wire net_3241;
wire net_2883;
wire net_2302;
wire net_998;
wire net_563;
wire net_2157;
wire net_1147;
wire net_3422;
wire net_2555;
wire net_199;
wire net_2789;
wire net_2681;
wire net_3027;
wire net_431;
wire net_2405;
wire net_2158;
wire net_835;
wire net_1687;
wire net_1762;
wire net_1181;
wire net_1266;
wire net_2368;
wire net_1452;
wire net_638;
wire net_1357;
wire net_2773;
wire net_2428;
wire net_909;
wire x793;
wire net_222;
wire net_313;
wire net_152;
wire net_932;
wire net_3105;
wire net_2895;
wire x279;
wire net_1788;
wire net_1243;
wire net_1660;
wire net_2138;
wire net_1484;
wire net_607;
wire net_258;
wire net_2477;
wire net_1783;
wire net_2935;
wire net_419;
wire net_1045;
wire net_2446;
wire net_1874;
wire net_1635;
wire net_972;
wire net_585;
wire net_936;
wire net_819;
wire net_1438;
wire net_785;
wire net_374;
wire net_3002;
wire net_1143;
wire net_1987;
wire net_1489;
wire net_854;
wire net_788;
wire net_2619;
wire net_214;
wire net_249;
wire net_3141;
wire net_1088;
wire net_1670;
wire net_2221;
wire net_3265;
wire net_2801;
wire net_1349;
wire net_2392;
wire net_2079;
wire net_979;
wire net_706;
wire net_1731;
wire net_2932;
wire net_2052;
wire net_156;
wire net_2015;
wire net_2768;
wire x2183;
wire net_1264;
wire net_2565;
wire net_2632;
wire net_551;
wire x609;
wire net_1040;
wire net_2547;
wire net_332;
wire net_1745;
wire net_1679;
wire net_3101;
wire net_3089;
wire net_3148;
wire net_3037;
wire x223;
wire net_1229;
wire net_2118;
wire net_463;
wire net_656;
wire net_2295;
wire net_1536;
wire net_1817;
wire net_197;
wire net_2560;
wire x258;
wire net_766;
wire net_2907;
wire net_1498;
wire net_1153;
wire net_1381;
wire net_3014;
wire net_1887;
wire x1817;
wire net_202;
wire net_1199;
wire net_3312;
wire net_1756;
wire net_2243;
wire net_379;
wire net_2208;
wire net_1569;
wire net_2595;
wire net_1383;
wire net_2751;
wire net_918;
wire net_3113;
wire net_949;
wire net_3133;
wire net_450;
wire net_289;
wire net_3047;
wire net_2559;
wire net_2614;
wire net_1642;
wire net_2657;
wire net_1358;
wire net_1683;
wire net_2629;
wire net_2486;
wire net_978;
wire net_2524;
wire net_1313;
wire net_2251;
wire x429;
wire net_1129;
wire net_3331;
wire net_1056;
wire net_1224;
wire net_2296;
wire net_1698;
wire net_768;
wire net_955;
wire net_1017;
wire net_2585;
wire net_1206;
wire net_3385;
wire net_357;
wire net_2044;
wire net_1996;
wire net_960;
wire net_2181;
wire x876;
wire net_1029;
wire net_1166;
wire net_908;
wire net_1789;
wire net_801;
wire net_519;
wire net_2620;
wire net_412;
wire net_2581;
wire net_1718;
wire net_838;
wire net_3219;
wire net_2986;
wire net_3162;
wire net_2694;
wire net_1873;
wire net_3118;
wire net_2129;
wire net_2096;
wire net_2697;
wire net_453;
wire net_581;
wire net_2899;
wire net_2576;
wire net_3180;
wire net_2352;
wire net_1038;
wire net_1829;
wire net_3249;
wire net_658;
wire net_1204;
wire net_2342;
wire net_2263;
wire net_734;
wire net_2544;
wire net_2090;
wire net_2325;
wire net_662;
wire net_3214;
wire net_1986;
wire net_862;
wire net_2086;
wire net_951;
wire net_50;
wire net_3186;
wire net_806;
wire net_3398;
wire net_2277;
wire net_2307;
wire net_342;
wire net_975;
wire net_612;
wire net_738;
wire net_892;
wire net_946;
wire net_1176;
wire net_1150;
wire net_504;
wire net_2966;
wire net_2676;
wire net_1253;
wire net_2194;
wire net_2500;
wire net_1076;
wire net_1751;
wire net_2006;
wire net_3406;
wire x2269;
wire net_1331;
wire net_1537;
wire x363;
wire net_3153;
wire net_681;
wire net_2130;
wire net_3362;
wire net_1148;
wire net_3120;
wire net_2434;
wire net_2032;
wire net_1448;
wire net_2214;
wire net_392;
wire net_3338;
wire net_118;
wire net_2467;
wire net_2382;
wire net_146;
wire net_1561;
wire net_2452;
wire net_2728;
wire net_417;
wire net_122;
wire net_3269;
wire x1192;
wire net_1502;
wire net_1940;
wire net_3337;
wire net_428;
wire net_2662;
wire net_94;
wire net_246;
wire x921;
wire net_1186;
wire x2242;
wire net_640;
wire net_482;
wire net_2888;
wire net_2216;
wire net_991;
wire net_3258;
wire x1280;
wire net_775;
wire net_149;
wire net_1378;
wire net_752;
wire net_3088;
wire net_387;
wire net_1773;
wire net_1473;
wire net_1600;
wire net_3275;
wire net_2531;
wire net_535;
wire net_498;
wire net_888;
wire net_2979;
wire net_676;
wire net_2772;
wire net_41;
wire net_1893;
wire net_1932;
wire net_1674;
wire net_1651;
wire net_2721;
wire net_577;
wire net_3401;
wire net_2375;
wire net_2637;
wire net_2538;
wire net_1023;
wire net_1806;
wire net_3234;
wire net_2550;
wire net_2447;
wire net_797;
wire net_2347;
wire net_301;
wire net_1957;
wire net_2360;
wire net_299;
wire net_1363;
wire net_1799;
wire net_1343;
wire net_2285;
wire net_1869;
wire net_2684;
wire net_2572;
wire net_2462;
wire net_182;
wire net_521;
wire net_60;
wire net_2414;
wire net_2754;
wire net_590;
wire net_337;
wire net_267;
wire net_2024;
wire net_1585;
wire net_1846;
wire net_3240;
wire net_3324;
wire x1222;
wire net_3254;
wire net_690;
wire net_523;
wire net_1370;
wire net_1435;
wire net_3260;
wire x1851;
wire net_407;
wire net_3207;
wire net_1736;
wire net_2204;
wire net_2716;
wire net_2371;
wire net_3375;
wire net_2492;
wire x1826;
wire net_2312;
wire net_1970;
wire net_1306;
wire net_351;
wire net_1669;
wire net_1858;
wire x1785;
wire net_2073;
wire net_1041;
wire net_3038;
wire net_2690;
wire net_2950;
wire net_1388;
wire net_2842;
wire net_791;
wire net_3158;
wire net_2828;
wire net_1257;
wire net_3239;
wire net_1419;
wire net_939;
wire net_2188;
wire net_824;
wire net_1051;
wire x1742;
wire net_3391;
wire net_2364;
wire net_1822;
wire net_2730;
wire net_942;
wire net_1631;
wire net_1337;
wire net_1182;
wire net_1624;
wire net_2791;
wire net_1981;
wire net_1972;
wire x780;
wire net_1515;
wire net_1218;
wire net_1638;
wire net_1950;
wire net_1573;
wire net_3126;
wire net_993;
wire net_1494;
wire net_3286;
wire net_361;
wire net_2890;
wire net_2154;
wire net_2421;
wire net_27;
wire x497;
wire net_1726;
wire net_317;
wire net_305;
wire net_856;
wire net_880;
wire net_1100;
wire net_1905;
wire net_1402;
wire net_3298;
wire net_3099;
wire net_2540;
wire net_1398;
wire net_2153;
wire net_1939;
wire net_2230;
wire net_1125;
wire net_2817;
wire net_3098;
wire net_144;
wire net_227;
wire net_2026;
wire x651;
wire net_1144;
wire net_1794;
wire net_2901;
wire net_162;
wire net_653;
wire net_1326;
wire net_3033;
wire net_134;
wire net_1022;
wire net_546;
wire x914;
wire net_1415;
wire net_2865;
wire net_2260;
wire net_3373;
wire net_3052;
wire net_2672;
wire net_3317;
wire net_3145;
wire net_2886;
wire net_1921;
wire net_702;
wire net_588;
wire net_3195;
wire net_1477;
wire net_3210;
wire x972;
wire net_3318;
wire net_2200;
wire net_2135;
wire net_1230;
wire net_667;
wire net_1157;
wire net_853;
wire net_236;
wire net_487;
wire net_212;
wire net_552;
wire net_914;
wire net_1787;
wire net_1542;
wire net_1172;
wire net_756;
wire net_1193;
wire net_1425;
wire net_875;
wire net_1122;
wire net_104;
wire net_1065;
wire net_2237;
wire net_3416;
wire net_72;
wire net_1813;
wire x1889;
wire net_2566;
wire net_1092;
wire net_627;
wire net_3100;
wire net_241;
wire net_917;
wire net_2039;
wire x316;
wire net_2874;
wire net_983;
wire net_355;
wire net_711;
wire net_599;
wire net_2225;
wire net_2993;
wire net_723;
wire net_1456;
wire net_3067;
wire x1312;
wire net_2483;
wire net_2227;
wire net_3111;
wire net_323;
wire net_2473;
wire net_963;
wire net_846;
wire net_3017;
wire x1343;
wire net_275;
wire net_399;
wire net_2914;
wire net_153;
wire net_2389;
wire net_1390;
wire net_218;
wire net_174;
wire net_2590;
wire net_2607;
wire net_1112;
wire net_3283;
wire net_1273;
wire net_562;
wire net_375;
wire net_364;
wire net_1137;
wire net_2506;
wire net_2114;
wire net_3172;
wire net_1831;
wire net_1482;
wire net_79;
wire net_3291;
wire net_3230;
wire net_2168;
wire net_3306;
wire net_2928;
wire net_2849;
wire x2049;
wire net_1885;
wire net_1030;
wire net_1485;
wire net_285;
wire net_3245;
wire net_1310;
wire net_2499;
wire net_254;
wire net_3171;
wire x208;
wire net_1297;
wire net_1501;
wire net_3003;
wire net_1304;
wire net_574;
wire net_2177;
wire x1405;
wire net_3357;
wire net_1247;
wire net_1969;
wire net_745;

// Start cells
INV_X8 inst_1783 ( .ZN(net_1611), .A(net_1610) );
NAND3_X2 inst_696 ( .ZN(net_2720), .A3(net_2719), .A2(net_2717), .A1(net_1880) );
CLKBUF_X2 inst_3311 ( .A(net_3268), .Z(net_3269) );
NAND2_X2 inst_1175 ( .ZN(net_101), .A1(net_86), .A2(x1047) );
NOR2_X2 inst_481 ( .ZN(net_2545), .A1(net_2544), .A2(net_2362) );
INV_X8 inst_1751 ( .ZN(net_130), .A(net_86) );
INV_X2 inst_2235 ( .ZN(net_294), .A(net_293) );
NAND2_X4 inst_779 ( .A2(net_1592), .ZN(net_1062), .A1(net_1061) );
NOR2_X2 inst_395 ( .A2(net_2603), .ZN(net_996), .A1(net_995) );
NAND2_X4 inst_841 ( .A1(net_2500), .ZN(net_1597), .A2(net_1596) );
INV_X2 inst_2205 ( .A(net_1864), .ZN(net_489) );
CLKBUF_X2 inst_2858 ( .A(net_2815), .Z(net_2816) );
NOR2_X2 inst_452 ( .ZN(net_1996), .A2(net_1994), .A1(net_453) );
NAND3_X2 inst_689 ( .ZN(net_2646), .A1(net_1835), .A2(net_1834), .A3(net_871) );
INV_X2 inst_2363 ( .A(net_2352), .ZN(net_1721) );
NOR2_X4 inst_214 ( .A2(net_2562), .A1(net_2129), .ZN(net_405) );
NAND2_X2 inst_1629 ( .ZN(net_2509), .A2(net_2507), .A1(net_1015) );
CLKBUF_X2 inst_3061 ( .A(net_3018), .Z(net_3019) );
NAND2_X2 inst_1558 ( .ZN(net_2115), .A1(net_1877), .A2(net_221) );
NAND4_X2 inst_548 ( .ZN(net_2331), .A1(net_1294), .A4(net_790), .A3(net_789), .A2(net_786) );
CLKBUF_X2 inst_2906 ( .A(net_2856), .Z(net_2864) );
NAND2_X4 inst_728 ( .A2(net_1494), .ZN(net_132), .A1(net_130) );
CLKBUF_X2 inst_3424 ( .A(net_3381), .Z(net_3382) );
CLKBUF_X2 inst_3121 ( .A(net_3058), .Z(net_3079) );
AOI21_X4 inst_2780 ( .ZN(net_2377), .B2(net_2376), .B1(net_2375), .A(net_2374) );
DFFR_X2 inst_2485 ( .D(net_1657), .Q(net_1504), .CK(net_2889), .RN(x2480) );
NAND2_X2 inst_1615 ( .ZN(net_2422), .A2(net_2160), .A1(net_1047) );
INV_X2 inst_2217 ( .ZN(net_545), .A(net_385) );
DFFR_X1 inst_2580 ( .D(net_2778), .CK(net_3367), .RN(x2480), .Q(x245) );
INV_X2 inst_2394 ( .A(net_2443), .ZN(net_2442) );
INV_X4 inst_2145 ( .A(net_2587), .ZN(net_2268) );
NAND2_X4 inst_850 ( .ZN(net_1662), .A2(net_1661), .A1(net_1340) );
NAND2_X4 inst_709 ( .A2(net_2111), .ZN(net_472), .A1(net_349) );
INV_X2 inst_2375 ( .ZN(net_1827), .A(x621) );
CLKBUF_X2 inst_3347 ( .A(net_2962), .Z(net_3305) );
CLKBUF_X2 inst_3130 ( .A(net_2855), .Z(net_3088) );
AND2_X2 inst_2844 ( .ZN(net_1125), .A1(net_1117), .A2(net_199) );
DFFR_X2 inst_2492 ( .D(net_2497), .Q(net_1480), .CK(net_2963), .RN(x2480) );
NAND2_X4 inst_920 ( .ZN(net_2033), .A1(net_1836), .A2(net_249) );
CLKBUF_X2 inst_3454 ( .A(net_3163), .Z(net_3412) );
INV_X4 inst_2054 ( .ZN(net_1301), .A(net_1300) );
NAND2_X2 inst_1228 ( .A1(net_1585), .A2(net_1473), .ZN(net_644) );
NAND2_X2 inst_1259 ( .A1(net_1942), .ZN(net_737), .A2(net_736) );
NAND4_X2 inst_521 ( .ZN(net_1151), .A1(net_1149), .A4(net_1135), .A3(net_1134), .A2(net_1133) );
INV_X8 inst_1796 ( .ZN(net_1904), .A(net_803) );
NAND2_X1 inst_1685 ( .ZN(net_496), .A1(net_495), .A2(net_348) );
DFFR_X2 inst_2511 ( .D(net_2228), .Q(net_1489), .CK(net_3290), .RN(x2480) );
INV_X16 inst_2438 ( .ZN(net_2408), .A(net_2407) );
NAND2_X2 inst_1655 ( .ZN(net_2619), .A1(net_2618), .A2(net_850) );
CLKBUF_X2 inst_2889 ( .A(net_2846), .Z(net_2847) );
NAND4_X2 inst_535 ( .ZN(net_1788), .A1(net_1787), .A2(net_1234), .A3(net_1136), .A4(net_603) );
AOI21_X4 inst_2772 ( .ZN(net_1614), .A(net_1613), .B2(net_1246), .B1(net_518) );
DFFR_X1 inst_2543 ( .QN(net_2801), .Q(net_1502), .D(net_943), .CK(net_3065), .RN(x2480) );
NOR2_X4 inst_237 ( .A1(net_2253), .A2(net_1322), .ZN(net_1106) );
NAND2_X2 inst_1670 ( .ZN(net_2703), .A2(net_2702), .A1(net_2699) );
INV_X4 inst_2189 ( .ZN(net_2662), .A(net_2658) );
NAND2_X4 inst_813 ( .A1(net_2296), .A2(net_1822), .ZN(net_1331) );
OAI21_X4 inst_51 ( .B1(net_1585), .A(net_650), .ZN(net_617), .B2(net_62) );
INV_X16 inst_2427 ( .ZN(net_2219), .A(net_2218) );
CLKBUF_X2 inst_2935 ( .A(net_2892), .Z(net_2893) );
NOR2_X4 inst_315 ( .ZN(net_2471), .A2(net_2470), .A1(net_917) );
INV_X8 inst_1837 ( .ZN(net_2470), .A(net_2469) );
NAND2_X2 inst_1066 ( .ZN(net_491), .A1(net_428), .A2(net_426) );
NAND2_X4 inst_974 ( .ZN(net_2353), .A2(net_2326), .A1(net_619) );
NOR2_X4 inst_216 ( .ZN(net_312), .A1(net_272), .A2(net_262) );
CLKBUF_X2 inst_3392 ( .A(net_3232), .Z(net_3350) );
CLKBUF_X2 inst_3317 ( .A(net_3274), .Z(net_3275) );
CLKBUF_X2 inst_3369 ( .A(net_3326), .Z(net_3327) );
INV_X2 inst_2342 ( .ZN(net_1347), .A(net_540) );
CLKBUF_X2 inst_3113 ( .A(net_2918), .Z(net_3071) );
CLKBUF_X2 inst_3291 ( .A(net_3248), .Z(net_3249) );
INV_X2 inst_2294 ( .ZN(net_34), .A(x1546) );
INV_X4 inst_2060 ( .A(net_1602), .ZN(net_1365) );
NAND2_X2 inst_1617 ( .A2(net_2519), .ZN(net_2431), .A1(net_2430) );
OAI21_X2 inst_151 ( .ZN(net_1595), .B1(net_1594), .A(net_1153), .B2(net_993) );
OAI21_X4 inst_64 ( .B1(net_2383), .ZN(net_1066), .B2(net_1008), .A(net_219) );
CLKBUF_X2 inst_3168 ( .A(net_3125), .Z(net_3126) );
INV_X2 inst_2256 ( .A(net_645), .ZN(net_138) );
NAND2_X4 inst_1001 ( .ZN(net_2493), .A2(net_2481), .A1(net_1432) );
INV_X2 inst_2385 ( .ZN(net_2164), .A(net_2157) );
INV_X2 inst_2336 ( .ZN(net_1246), .A(net_1241) );
INV_X4 inst_2106 ( .ZN(net_1834), .A(net_275) );
NAND2_X4 inst_743 ( .A1(net_2320), .ZN(net_689), .A2(net_209) );
NOR2_X2 inst_415 ( .ZN(net_1265), .A2(net_1264), .A1(net_483) );
AOI22_X2 inst_2723 ( .A2(net_2768), .ZN(net_1145), .A1(net_295), .B1(net_126), .B2(x1466) );
CLKBUF_X2 inst_3033 ( .A(net_2990), .Z(net_2991) );
INV_X8 inst_1795 ( .ZN(net_1858), .A(net_1857) );
NAND2_X4 inst_828 ( .A2(net_2380), .ZN(net_1445), .A1(net_1431) );
CLKBUF_X2 inst_2925 ( .A(net_2854), .Z(net_2883) );
CLKBUF_X2 inst_3318 ( .A(net_3275), .Z(net_3276) );
NOR2_X4 inst_223 ( .A1(net_1651), .ZN(net_799), .A2(net_795) );
INV_X8 inst_1828 ( .ZN(net_2399), .A(net_2398) );
INV_X4 inst_2072 ( .ZN(net_1579), .A(net_1578) );
NAND2_X2 inst_1603 ( .ZN(net_2354), .A2(net_2323), .A1(net_1410) );
INV_X8 inst_1809 ( .A(net_2727), .ZN(net_2118) );
NOR2_X2 inst_340 ( .A2(net_2538), .A1(net_529), .ZN(net_453) );
CLKBUF_X2 inst_3388 ( .A(net_3001), .Z(net_3346) );
INV_X16 inst_2420 ( .A(net_2327), .ZN(net_1943) );
NAND2_X2 inst_1561 ( .A1(net_2320), .ZN(net_2124), .A2(net_173) );
OAI21_X2 inst_158 ( .B2(net_2351), .ZN(net_1900), .A(net_1862), .B1(net_861) );
OAI21_X2 inst_141 ( .ZN(net_1337), .A(net_1336), .B1(net_801), .B2(net_556) );
DFFR_X2 inst_2520 ( .D(net_2234), .Q(net_1505), .CK(net_2906), .RN(x2480) );
INV_X4 inst_2104 ( .A(net_1824), .ZN(net_1820) );
NAND2_X2 inst_1322 ( .A1(net_1437), .A2(net_1196), .ZN(net_970) );
DFFR_X1 inst_2573 ( .D(net_2779), .CK(net_3402), .RN(x2480), .Q(x302) );
NAND2_X2 inst_1490 ( .A1(net_2348), .ZN(net_1754), .A2(net_1753) );
NAND4_X4 inst_507 ( .ZN(net_2279), .A4(net_1945), .A3(net_1944), .A2(net_1940), .A1(net_1939) );
NAND3_X4 inst_571 ( .ZN(net_1762), .A1(net_311), .A2(net_269), .A3(net_253) );
INV_X4 inst_1974 ( .A(net_1588), .ZN(net_782) );
INV_X4 inst_2017 ( .ZN(net_1035), .A(net_1032) );
NAND2_X4 inst_884 ( .ZN(net_1842), .A2(net_766), .A1(net_765) );
NAND2_X2 inst_1154 ( .A2(net_1527), .ZN(net_128), .A1(net_117) );
NAND2_X4 inst_711 ( .A2(net_1582), .A1(net_655), .ZN(net_527) );
NAND2_X4 inst_827 ( .A1(net_2440), .A2(net_2426), .ZN(net_1438) );
INV_X4 inst_2096 ( .ZN(net_1764), .A(net_1763) );
NAND4_X2 inst_552 ( .ZN(net_2527), .A3(net_1669), .A1(net_1436), .A4(net_838), .A2(net_837) );
CLKBUF_X2 inst_3050 ( .A(net_3007), .Z(net_3008) );
NOR2_X2 inst_469 ( .ZN(net_2173), .A2(net_1608), .A1(net_441) );
CLKBUF_X2 inst_3040 ( .A(net_2997), .Z(net_2998) );
CLKBUF_X2 inst_3019 ( .A(net_2976), .Z(net_2977) );
CLKBUF_X2 inst_2980 ( .A(net_2937), .Z(net_2938) );
INV_X2 inst_2327 ( .A(net_1678), .ZN(net_1004) );
NAND2_X2 inst_1564 ( .A2(net_2204), .ZN(net_2139), .A1(net_833) );
OAI22_X4 inst_18 ( .B2(net_2807), .ZN(net_1828), .A2(net_1827), .B1(net_1826), .A1(net_1825) );
NAND2_X4 inst_915 ( .A1(net_2235), .A2(net_2233), .ZN(net_2016) );
INV_X4 inst_1941 ( .A(net_1589), .ZN(net_156) );
INV_X2 inst_2263 ( .ZN(net_64), .A(x1427) );
DFFR_X1 inst_2607 ( .D(net_2754), .CK(net_3397), .RN(x2480), .Q(x287) );
INV_X2 inst_2339 ( .A(net_2484), .ZN(net_1272) );
OR2_X2 inst_9 ( .A2(net_2795), .A1(net_1586), .ZN(net_859) );
OAI21_X2 inst_113 ( .A(net_724), .B2(net_319), .ZN(net_261), .B1(net_154) );
NOR2_X2 inst_356 ( .A1(net_2693), .A2(net_2157), .ZN(net_373) );
CLKBUF_X2 inst_3358 ( .A(net_3315), .Z(net_3316) );
NAND2_X2 inst_1216 ( .A1(net_1585), .A2(net_1485), .ZN(net_628) );
NAND2_X4 inst_952 ( .ZN(net_2229), .A1(net_2228), .A2(net_2225) );
NAND2_X2 inst_1668 ( .ZN(net_2696), .A1(net_2695), .A2(net_2135) );
NAND2_X2 inst_1594 ( .ZN(net_2306), .A2(net_2305), .A1(net_2304) );
NAND2_X4 inst_721 ( .A1(net_625), .ZN(net_245), .A2(net_97) );
NAND2_X4 inst_902 ( .ZN(net_1949), .A2(net_1938), .A1(net_1936) );
NOR2_X4 inst_293 ( .A1(net_2727), .ZN(net_2135), .A2(net_1021) );
NAND2_X4 inst_778 ( .A1(net_2259), .A2(net_1541), .ZN(net_1050) );
CLKBUF_X2 inst_3009 ( .A(net_2966), .Z(net_2967) );
NAND2_X2 inst_1366 ( .A2(net_1203), .ZN(net_1170), .A1(net_898) );
NAND2_X2 inst_1544 ( .ZN(net_2060), .A1(net_2058), .A2(net_1014) );
INV_X4 inst_1935 ( .A(net_1076), .ZN(net_142) );
CLKBUF_X2 inst_3102 ( .A(net_3059), .Z(net_3060) );
AOI22_X4 inst_2695 ( .ZN(net_1803), .B1(net_985), .A2(net_756), .A1(net_755), .B2(net_718) );
INV_X4 inst_1915 ( .ZN(net_279), .A(net_278) );
AOI21_X2 inst_2794 ( .B2(net_2538), .B1(net_2457), .ZN(net_876), .A(net_875) );
DFFR_X1 inst_2625 ( .Q(net_2775), .D(net_182), .CK(net_3297), .RN(x2480) );
INV_X4 inst_2063 ( .ZN(net_1431), .A(net_1430) );
NAND2_X2 inst_1254 ( .ZN(net_726), .A2(net_721), .A1(net_631) );
CLKBUF_X2 inst_3148 ( .A(net_3105), .Z(net_3106) );
CLKBUF_X2 inst_2953 ( .A(net_2910), .Z(net_2911) );
INV_X4 inst_2140 ( .ZN(net_2186), .A(net_2183) );
CLKBUF_X2 inst_3329 ( .A(net_3286), .Z(net_3287) );
NAND2_X4 inst_781 ( .A1(net_2196), .A2(net_2194), .ZN(net_1073) );
INV_X8 inst_1811 ( .ZN(net_2133), .A(net_2132) );
OAI21_X4 inst_98 ( .ZN(net_2348), .B2(net_2347), .B1(net_2345), .A(net_2344) );
CLKBUF_X2 inst_3440 ( .A(net_3395), .Z(net_3398) );
CLKBUF_X2 inst_3087 ( .A(net_3044), .Z(net_3045) );
INV_X4 inst_2036 ( .ZN(net_1180), .A(net_1179) );
CLKBUF_X2 inst_3026 ( .A(net_2983), .Z(net_2984) );
NAND2_X4 inst_959 ( .A2(net_2587), .ZN(net_2271), .A1(net_867) );
AND2_X2 inst_2847 ( .A1(net_2303), .ZN(net_1206), .A2(net_298) );
NAND2_X2 inst_1442 ( .A2(net_2023), .A1(net_2001), .ZN(net_1462) );
NOR2_X4 inst_332 ( .ZN(net_2705), .A1(net_2704), .A2(net_967) );
INV_X4 inst_2049 ( .ZN(net_1275), .A(net_1274) );
NAND2_X4 inst_868 ( .ZN(net_1746), .A2(net_1745), .A1(net_1744) );
OAI21_X2 inst_163 ( .B2(net_2784), .ZN(net_2107), .A(net_2003), .B1(net_169) );
NOR2_X2 inst_394 ( .A2(net_2693), .A1(net_2425), .ZN(net_967) );
INV_X4 inst_2132 ( .ZN(net_2094), .A(net_2093) );
NAND2_X2 inst_1289 ( .ZN(net_2147), .A2(net_1959), .A1(net_334) );
INV_X4 inst_1928 ( .ZN(net_295), .A(net_126) );
NAND2_X2 inst_1559 ( .ZN(net_2116), .A1(net_247), .A2(net_158) );
INV_X4 inst_1967 ( .A(net_1672), .ZN(net_746) );
NOR3_X2 inst_201 ( .A2(net_2433), .A1(net_1889), .A3(net_1428), .ZN(net_392) );
NAND2_X4 inst_927 ( .ZN(net_2088), .A2(net_2087), .A1(net_945) );
NAND3_X2 inst_605 ( .A1(net_2165), .A2(net_1850), .ZN(net_958), .A3(net_957) );
NAND2_X2 inst_1084 ( .A1(net_2402), .A2(net_2336), .ZN(net_434) );
NOR2_X4 inst_304 ( .A2(net_2684), .A1(net_2683), .ZN(net_2283) );
INV_X8 inst_1814 ( .ZN(net_2165), .A(net_2157) );
CLKBUF_X2 inst_3245 ( .A(net_3077), .Z(net_3203) );
AOI21_X2 inst_2799 ( .A(net_2433), .B2(net_1286), .ZN(net_1039), .B1(net_519) );
NAND2_X4 inst_752 ( .A2(net_1127), .ZN(net_752), .A1(net_696) );
CLKBUF_X2 inst_3202 ( .A(net_3159), .Z(net_3160) );
INV_X4 inst_1947 ( .A(net_873), .ZN(net_81) );
NAND2_X1 inst_1719 ( .A1(net_1808), .A2(net_1805), .ZN(net_1319) );
NAND2_X2 inst_1488 ( .ZN(net_1749), .A2(net_1748), .A1(net_1747) );
NAND2_X4 inst_1027 ( .ZN(net_2675), .A2(net_2674), .A1(net_2673) );
OAI21_X4 inst_73 ( .ZN(net_1424), .B2(net_1421), .B1(net_1245), .A(net_884) );
NAND2_X2 inst_1143 ( .A1(net_246), .A2(net_187), .ZN(net_184) );
INV_X4 inst_1951 ( .A(net_760), .ZN(net_593) );
NAND2_X2 inst_1345 ( .A2(net_1666), .ZN(net_1070), .A1(net_1069) );
NOR2_X2 inst_378 ( .A1(net_1730), .A2(net_1407), .ZN(net_808) );
NAND2_X2 inst_1384 ( .ZN(net_1256), .A1(net_841), .A2(net_681) );
CLKBUF_X2 inst_2947 ( .A(net_2904), .Z(net_2905) );
INV_X4 inst_2118 ( .ZN(net_1959), .A(net_1958) );
INV_X4 inst_2048 ( .ZN(net_1269), .A(net_1268) );
NAND2_X4 inst_890 ( .A2(net_2269), .ZN(net_1870), .A1(net_661) );
INV_X32 inst_2200 ( .ZN(net_2237), .A(net_2236) );
CLKBUF_X2 inst_2948 ( .A(net_2905), .Z(net_2906) );
INV_X4 inst_1851 ( .A(net_1180), .ZN(net_538) );
NOR2_X2 inst_361 ( .ZN(net_238), .A2(net_237), .A1(net_229) );
NAND2_X2 inst_1168 ( .ZN(net_691), .A1(net_86), .A2(x663) );
CLKBUF_X2 inst_3400 ( .A(net_3357), .Z(net_3358) );
NAND2_X4 inst_1016 ( .ZN(net_2584), .A2(net_1093), .A1(net_888) );
NAND2_X2 inst_1538 ( .A2(net_2387), .ZN(net_2007), .A1(net_2006) );
NAND3_X2 inst_659 ( .A2(net_2267), .A3(net_2062), .ZN(net_2053), .A1(net_607) );
NOR2_X4 inst_250 ( .A1(net_2076), .A2(net_1654), .ZN(net_1241) );
NAND2_X4 inst_848 ( .ZN(net_1638), .A2(net_1509), .A1(net_980) );
INV_X4 inst_1931 ( .A(net_2237), .ZN(net_240) );
CLKBUF_X2 inst_3002 ( .A(net_2959), .Z(net_2960) );
DFFR_X2 inst_2479 ( .D(net_1554), .Q(net_1494), .CK(net_3130), .RN(x2480) );
INV_X4 inst_2179 ( .ZN(net_2548), .A(net_2547) );
DFFR_X1 inst_2578 ( .D(net_2773), .CK(net_2852), .RN(x2480), .Q(x439) );
NAND2_X4 inst_786 ( .A1(net_1258), .ZN(net_1096), .A2(x921) );
CLKBUF_X2 inst_3362 ( .A(net_3319), .Z(net_3320) );
NAND2_X2 inst_1161 ( .A1(net_133), .ZN(net_119), .A2(net_71) );
DFFR_X1 inst_2539 ( .D(net_1150), .Q(net_79), .CK(net_3086), .RN(x2480) );
NAND2_X2 inst_1523 ( .ZN(net_1952), .A2(net_1951), .A1(net_1950) );
CLKBUF_X2 inst_2940 ( .A(net_2817), .Z(net_2898) );
INV_X4 inst_1996 ( .A(net_2227), .ZN(net_908) );
NAND2_X2 inst_1554 ( .A1(net_2458), .ZN(net_2101), .A2(net_179) );
NAND2_X2 inst_1542 ( .A2(net_2061), .ZN(net_2041), .A1(net_2004) );
NAND2_X2 inst_1048 ( .A2(net_2137), .ZN(net_553), .A1(net_537) );
CLKBUF_X2 inst_3199 ( .A(net_3156), .Z(net_3157) );
AOI21_X2 inst_2797 ( .B2(net_1816), .A(net_1137), .ZN(net_1029), .B1(net_683) );
XNOR2_X2 inst_2 ( .ZN(net_2063), .B(net_1514), .A(net_712) );
CLKBUF_X2 inst_3340 ( .A(net_2940), .Z(net_3298) );
NAND3_X2 inst_644 ( .ZN(net_1798), .A1(net_1797), .A3(net_974), .A2(net_973) );
CLKBUF_X2 inst_3431 ( .A(net_3388), .Z(net_3389) );
NAND2_X2 inst_1581 ( .A2(net_2295), .ZN(net_2216), .A1(net_1822) );
INV_X2 inst_2270 ( .ZN(net_57), .A(x1980) );
INV_X2 inst_2388 ( .ZN(net_2225), .A(net_2224) );
INV_X4 inst_2085 ( .A(net_1666), .ZN(net_1654) );
INV_X2 inst_2401 ( .ZN(net_2573), .A(net_2572) );
NAND2_X2 inst_1380 ( .A2(net_2318), .ZN(net_1235), .A1(net_1007) );
AOI21_X2 inst_2806 ( .A(net_1567), .ZN(net_1285), .B1(net_1281), .B2(net_673) );
INV_X2 inst_2312 ( .ZN(net_798), .A(net_794) );
NAND3_X4 inst_578 ( .ZN(net_2258), .A1(net_2256), .A3(net_614), .A2(net_613) );
NAND2_X4 inst_888 ( .A2(net_2326), .ZN(net_1861), .A1(net_927) );
INV_X8 inst_1769 ( .A(net_2054), .ZN(net_1083) );
DFFR_X1 inst_2634 ( .D(net_71), .CK(net_3194), .RN(x2480), .Q(x49) );
INV_X2 inst_2241 ( .A(net_1942), .ZN(net_193) );
INV_X4 inst_2182 ( .ZN(net_2608), .A(net_2370) );
DFFR_X1 inst_2581 ( .D(net_2761), .CK(net_3334), .RN(x2480), .Q(x216) );
NAND4_X2 inst_556 ( .ZN(net_2640), .A2(net_2639), .A1(net_1397), .A4(net_1337), .A3(net_901) );
NAND3_X2 inst_650 ( .A2(net_2316), .A1(net_2315), .ZN(net_1938), .A3(net_1937) );
NOR2_X4 inst_289 ( .A1(net_2592), .ZN(net_2084), .A2(net_159) );
INV_X4 inst_2164 ( .A(net_2805), .ZN(net_2418) );
NAND2_X4 inst_987 ( .ZN(net_2403), .A1(net_1989), .A2(net_1038) );
NAND2_X2 inst_1498 ( .A1(net_2696), .A2(net_2290), .ZN(net_1800) );
NOR2_X2 inst_432 ( .ZN(net_1443), .A2(net_1442), .A1(net_1441) );
NAND3_X2 inst_679 ( .ZN(net_2456), .A1(net_2455), .A3(net_1638), .A2(net_1164) );
NOR2_X2 inst_420 ( .A2(net_2416), .ZN(net_1348), .A1(net_1016) );
NOR2_X4 inst_282 ( .ZN(net_1869), .A2(net_1868), .A1(net_1553) );
NAND2_X2 inst_1358 ( .ZN(net_1131), .A2(net_721), .A1(net_664) );
CLKBUF_X2 inst_3006 ( .A(net_2860), .Z(net_2964) );
CLKBUF_X2 inst_3265 ( .A(net_3222), .Z(net_3223) );
INV_X2 inst_2322 ( .ZN(net_931), .A(net_930) );
NAND4_X2 inst_513 ( .A2(net_2397), .ZN(net_889), .A4(net_414), .A1(net_370), .A3(net_351) );
CLKBUF_X2 inst_3364 ( .A(net_3254), .Z(net_3322) );
CLKBUF_X2 inst_3266 ( .A(net_3223), .Z(net_3224) );
CLKBUF_X2 inst_3171 ( .A(net_3128), .Z(net_3129) );
NAND2_X2 inst_1351 ( .A2(net_2386), .A1(net_2321), .ZN(net_1097) );
OAI221_X1 inst_44 ( .B2(net_2031), .B1(net_327), .ZN(net_325), .C2(net_319), .A(net_303), .C1(net_171) );
CLKBUF_X2 inst_3300 ( .A(net_3257), .Z(net_3258) );
NAND2_X2 inst_1630 ( .ZN(net_2511), .A1(net_1446), .A2(net_1073) );
NAND2_X2 inst_1305 ( .A2(net_1547), .ZN(net_914), .A1(net_395) );
NOR2_X2 inst_371 ( .A1(net_2567), .A2(net_2396), .ZN(net_768) );
NAND2_X2 inst_1586 ( .ZN(net_2255), .A1(net_2254), .A2(net_1415) );
NOR2_X4 inst_314 ( .A2(net_2516), .ZN(net_2464), .A1(net_343) );
CLKBUF_X2 inst_3385 ( .A(net_3342), .Z(net_3343) );
CLKBUF_X2 inst_3225 ( .A(net_3182), .Z(net_3183) );
CLKBUF_X2 inst_3182 ( .A(net_3139), .Z(net_3140) );
NOR2_X2 inst_435 ( .A2(net_2179), .ZN(net_1582), .A1(net_849) );
NAND2_X2 inst_1572 ( .ZN(net_2174), .A2(net_2173), .A1(net_2172) );
NAND3_X2 inst_597 ( .A3(net_2071), .A1(net_1654), .ZN(net_840), .A2(net_361) );
CLKBUF_X2 inst_2866 ( .A(net_2823), .Z(net_2824) );
NAND2_X4 inst_774 ( .A2(net_1853), .ZN(net_1027), .A1(net_1026) );
CLKBUF_X2 inst_3307 ( .A(net_3264), .Z(net_3265) );
INV_X2 inst_2292 ( .ZN(net_36), .A(x850) );
NAND2_X2 inst_1587 ( .A2(net_2323), .ZN(net_2263), .A1(net_2262) );
NAND2_X2 inst_1185 ( .ZN(net_1212), .A1(net_98), .A2(x1126) );
NAND2_X4 inst_838 ( .A1(net_2259), .ZN(net_1576), .A2(net_1519) );
NAND3_X2 inst_628 ( .A3(net_2005), .A2(net_1687), .ZN(net_1562), .A1(net_1561) );
CLKBUF_X2 inst_3013 ( .A(net_2845), .Z(net_2971) );
AOI22_X2 inst_2748 ( .ZN(net_2604), .A2(net_1547), .B1(net_1291), .B2(net_1290), .A1(net_1289) );
INV_X4 inst_1923 ( .A(net_1845), .ZN(net_178) );
NOR2_X2 inst_472 ( .A1(net_2726), .ZN(net_2358), .A2(net_2357) );
NOR2_X2 inst_447 ( .A2(net_1974), .A1(net_1965), .ZN(net_1801) );
NOR2_X2 inst_457 ( .A2(net_2365), .ZN(net_2037), .A1(net_1028) );
AOI21_X4 inst_2766 ( .B2(net_2563), .B1(net_2462), .A(net_2099), .ZN(net_1095) );
INV_X8 inst_1738 ( .ZN(net_350), .A(net_338) );
NAND2_X2 inst_1508 ( .ZN(net_1853), .A2(net_1852), .A1(net_1703) );
AOI21_X2 inst_2802 ( .B1(net_1964), .B2(net_1280), .ZN(net_1202), .A(net_392) );
DFFR_X1 inst_2623 ( .Q(net_2765), .D(net_1757), .CK(net_3009), .RN(x2480) );
CLKBUF_X2 inst_3092 ( .A(net_3049), .Z(net_3050) );
NAND2_X2 inst_1391 ( .A2(net_2409), .ZN(net_1279), .A1(net_1156) );
NAND2_X2 inst_1222 ( .A1(net_1585), .A2(net_1543), .ZN(net_638) );
NAND3_X2 inst_665 ( .A3(net_2682), .A1(net_2681), .ZN(net_2209), .A2(net_2037) );
NAND2_X2 inst_1405 ( .ZN(net_1328), .A2(net_1327), .A1(net_1325) );
CLKBUF_X2 inst_3407 ( .A(net_3364), .Z(net_3365) );
AOI22_X2 inst_2734 ( .A2(net_2320), .ZN(net_2006), .A1(net_1098), .B1(net_1051), .B2(net_242) );
NAND2_X2 inst_1073 ( .A1(net_991), .A2(net_707), .ZN(net_476) );
INV_X2 inst_2323 ( .ZN(net_933), .A(net_930) );
CLKBUF_X2 inst_3395 ( .A(net_3352), .Z(net_3353) );
NAND2_X2 inst_1130 ( .A2(net_2237), .ZN(net_204), .A1(net_203) );
AOI22_X2 inst_2749 ( .ZN(net_2745), .A2(net_1943), .B2(net_217), .A1(net_216), .B1(net_163) );
NAND2_X2 inst_1449 ( .A1(net_1567), .ZN(net_1565), .A2(net_382) );
OAI21_X2 inst_127 ( .ZN(net_877), .A(net_529), .B2(net_488), .B1(net_484) );
NAND2_X4 inst_855 ( .ZN(net_1675), .A2(net_1674), .A1(net_1673) );
INV_X4 inst_2039 ( .A(net_2078), .ZN(net_1200) );
OAI21_X2 inst_146 ( .B1(net_1682), .B2(net_1414), .ZN(net_1408), .A(net_364) );
CLKBUF_X2 inst_3233 ( .A(net_3041), .Z(net_3191) );
INV_X4 inst_2013 ( .ZN(net_1014), .A(net_1012) );
OAI211_X2 inst_187 ( .C1(net_2493), .B(net_2206), .A(net_2011), .ZN(net_1030), .C2(net_915) );
NOR3_X2 inst_206 ( .ZN(net_1396), .A3(net_1395), .A2(net_1393), .A1(net_1347) );
CLKBUF_X2 inst_3029 ( .A(net_2986), .Z(net_2987) );
NAND2_X2 inst_1268 ( .A2(net_1163), .ZN(net_771), .A1(net_444) );
OAI21_X2 inst_122 ( .B1(net_2383), .B2(net_1690), .A(net_1381), .ZN(net_760) );
AOI222_X1 inst_2756 ( .B2(net_2321), .A2(net_1410), .C2(net_736), .B1(net_721), .ZN(net_676), .C1(net_619), .A1(net_158) );
NAND2_X2 inst_1196 ( .A1(net_2239), .ZN(net_582), .A2(net_252) );
NOR2_X2 inst_405 ( .ZN(net_1124), .A2(net_1123), .A1(net_1122) );
NAND2_X1 inst_1731 ( .ZN(net_2737), .A1(net_2736), .A2(net_716) );
NOR2_X1 inst_492 ( .A1(net_2537), .A2(net_1509), .ZN(net_863) );
NAND2_X4 inst_817 ( .A1(net_1752), .ZN(net_1374), .A2(net_280) );
NOR2_X4 inst_326 ( .ZN(net_2621), .A1(net_1607), .A2(net_371) );
CLKBUF_X2 inst_3428 ( .A(net_3029), .Z(net_3386) );
INV_X4 inst_2194 ( .ZN(net_2700), .A(net_2697) );
NAND2_X2 inst_1363 ( .A1(net_2118), .ZN(net_1154), .A2(net_780) );
NAND4_X2 inst_518 ( .A3(net_1696), .A4(net_1121), .A2(net_1100), .ZN(net_1093), .A1(net_1067) );
CLKBUF_X2 inst_3336 ( .A(net_3293), .Z(net_3294) );
CLKBUF_X2 inst_2960 ( .A(net_2917), .Z(net_2918) );
INV_X4 inst_1909 ( .ZN(net_271), .A(net_263) );
CLKBUF_X2 inst_3293 ( .A(net_3250), .Z(net_3251) );
INV_X2 inst_2306 ( .ZN(net_756), .A(net_720) );
AND2_X4 inst_2837 ( .ZN(net_2355), .A2(net_2354), .A1(net_2353) );
INV_X2 inst_2345 ( .ZN(net_1417), .A(net_1411) );
OAI21_X4 inst_82 ( .ZN(net_1877), .A(net_638), .B2(net_117), .B1(net_30) );
NAND2_X2 inst_1646 ( .ZN(net_2591), .A2(net_2589), .A1(net_2386) );
INV_X8 inst_1845 ( .ZN(net_2567), .A(net_2557) );
OAI21_X2 inst_108 ( .A(net_799), .B1(net_798), .ZN(net_543), .B2(net_473) );
INV_X4 inst_2176 ( .ZN(net_2512), .A(net_2511) );
CLKBUF_X2 inst_2892 ( .A(net_2849), .Z(net_2850) );
NAND2_X2 inst_1121 ( .A2(net_1943), .A1(net_1051), .ZN(net_219) );
NAND2_X2 inst_1102 ( .A1(net_2685), .A2(net_670), .ZN(net_335) );
CLKBUF_X2 inst_3161 ( .A(net_3118), .Z(net_3119) );
CLKBUF_X2 inst_3187 ( .A(net_3144), .Z(net_3145) );
NAND2_X2 inst_1354 ( .A1(net_2738), .A2(net_2524), .ZN(net_1114) );
NAND2_X2 inst_1429 ( .A2(net_2488), .ZN(net_1385), .A1(net_1040) );
NAND2_X4 inst_970 ( .ZN(net_2340), .A1(net_411), .A2(net_372) );
NOR2_X4 inst_307 ( .ZN(net_2301), .A2(net_2092), .A1(net_2091) );
NAND2_X2 inst_1278 ( .A2(net_2237), .ZN(net_827), .A1(net_136) );
NAND3_X2 inst_638 ( .ZN(net_1677), .A3(net_1674), .A1(net_1673), .A2(net_1588) );
NAND2_X4 inst_749 ( .ZN(net_743), .A1(net_326), .A2(net_314) );
NAND3_X2 inst_586 ( .A3(net_2561), .A1(net_1934), .ZN(net_430), .A2(net_346) );
AOI21_X2 inst_2816 ( .ZN(net_2292), .B1(net_910), .B2(net_761), .A(net_549) );
NAND3_X1 inst_702 ( .A3(net_2219), .ZN(net_1433), .A1(net_1432), .A2(net_449) );
INV_X4 inst_2034 ( .A(net_1746), .ZN(net_1166) );
NAND2_X2 inst_1505 ( .ZN(net_1845), .A1(net_1844), .A2(net_859) );
NAND2_X4 inst_717 ( .A1(net_623), .ZN(net_244), .A2(net_99) );
NOR2_X4 inst_276 ( .ZN(net_1785), .A2(net_1784), .A1(net_465) );
DFFR_X2 inst_2482 ( .QN(net_2809), .D(net_572), .CK(net_2830), .RN(x2480) );
INV_X4 inst_2127 ( .ZN(net_2023), .A(net_2017) );
NAND2_X4 inst_1030 ( .ZN(net_2691), .A1(net_2690), .A2(net_2190) );
CLKBUF_X2 inst_2957 ( .A(net_2914), .Z(net_2915) );
DFFR_X1 inst_2649 ( .D(net_1536), .CK(net_3238), .RN(x2480), .Q(x136) );
DFFR_X1 inst_2591 ( .D(net_2768), .CK(net_3349), .RN(x2480), .Q(x144) );
CLKBUF_X2 inst_3275 ( .A(net_2921), .Z(net_3233) );
CLKBUF_X2 inst_3339 ( .A(net_3296), .Z(net_3297) );
NAND2_X2 inst_1466 ( .ZN(net_1655), .A1(net_1260), .A2(net_736) );
AND2_X2 inst_2841 ( .ZN(net_963), .A1(net_245), .A2(net_187) );
NAND2_X1 inst_1726 ( .A1(net_2399), .A2(net_1918), .ZN(net_1817) );
AOI22_X2 inst_2711 ( .A2(net_2761), .A1(net_295), .ZN(net_293), .B1(net_126), .B2(x1645) );
DFFR_X1 inst_2652 ( .D(net_1524), .CK(net_2840), .RN(x2480), .Q(x405) );
INV_X2 inst_2268 ( .ZN(net_59), .A(x1214) );
NAND2_X2 inst_1373 ( .A1(net_2366), .A2(net_1901), .ZN(net_1198) );
AOI222_X1 inst_2753 ( .C1(net_1943), .A2(net_736), .ZN(net_303), .C2(net_247), .B2(net_244), .B1(net_158), .A1(net_149) );
INV_X1 inst_2458 ( .A(net_1969), .ZN(net_677) );
NAND2_X2 inst_1203 ( .A1(net_2318), .A2(net_2239), .ZN(net_600) );
NAND2_X4 inst_802 ( .A1(net_1902), .ZN(net_1247), .A2(net_823) );
NOR2_X4 inst_296 ( .A2(net_2693), .ZN(net_2160), .A1(net_2159) );
OAI21_X4 inst_91 ( .ZN(net_2190), .B2(net_2189), .A(net_850), .B1(net_480) );
INV_X8 inst_1762 ( .A(net_2132), .ZN(net_736) );
NAND2_X4 inst_905 ( .ZN(net_1961), .A2(net_1788), .A1(net_1247) );
OAI21_X2 inst_132 ( .ZN(net_1058), .B2(net_1057), .A(net_799), .B1(net_604) );
INV_X4 inst_2023 ( .ZN(net_1086), .A(net_1081) );
CLKBUF_X2 inst_3155 ( .A(net_3112), .Z(net_3113) );
CLKBUF_X2 inst_3134 ( .A(net_2889), .Z(net_3092) );
AOI21_X4 inst_2779 ( .ZN(net_2291), .B2(net_2290), .B1(net_2289), .A(net_2285) );
NAND2_X4 inst_1006 ( .ZN(net_2523), .A1(net_1667), .A2(net_1271) );
INV_X4 inst_1985 ( .ZN(net_831), .A(net_830) );
NAND2_X1 inst_1703 ( .A1(net_632), .ZN(net_109), .A2(x1244) );
INV_X8 inst_1759 ( .A(net_1684), .ZN(net_686) );
CLKBUF_X2 inst_2928 ( .A(net_2827), .Z(net_2886) );
DFFR_X1 inst_2615 ( .Q(net_2753), .D(net_2107), .CK(net_3325), .RN(x2480) );
NOR2_X2 inst_400 ( .A2(net_2216), .A1(net_1723), .ZN(net_1041) );
CLKBUF_X2 inst_2991 ( .A(net_2948), .Z(net_2949) );
DFFR_X2 inst_2532 ( .QN(net_2802), .D(net_94), .CK(net_3181), .RN(x2480) );
CLKBUF_X2 inst_3463 ( .A(net_3257), .Z(net_3421) );
INV_X1 inst_2463 ( .A(net_1577), .ZN(net_1377) );
NAND3_X2 inst_614 ( .A2(net_2283), .A1(net_2203), .ZN(net_1255), .A3(net_677) );
INV_X4 inst_1896 ( .A(net_2408), .ZN(net_504) );
NOR2_X4 inst_261 ( .A2(net_2362), .A1(net_1720), .ZN(net_1452) );
NAND2_X2 inst_1464 ( .ZN(net_1637), .A2(net_1636), .A1(net_1634) );
NAND2_X2 inst_1247 ( .A1(net_2551), .A2(net_1820), .ZN(net_700) );
NAND2_X4 inst_1031 ( .ZN(net_2693), .A2(net_2692), .A1(net_2147) );
NAND2_X4 inst_945 ( .ZN(net_2182), .A1(net_2181), .A2(net_83) );
NOR2_X4 inst_268 ( .A2(net_2325), .ZN(net_1606), .A1(net_1365) );
NAND2_X2 inst_1518 ( .ZN(net_1935), .A2(net_1933), .A1(net_1407) );
NOR2_X2 inst_369 ( .A1(net_2138), .A2(net_1767), .ZN(net_710) );
INV_X4 inst_1900 ( .ZN(net_342), .A(net_340) );
NAND2_X2 inst_1493 ( .A1(net_2386), .ZN(net_1756), .A2(net_173) );
NOR2_X4 inst_327 ( .ZN(net_2629), .A2(net_2628), .A1(net_2081) );
NAND2_X2 inst_1308 ( .A1(net_1312), .ZN(net_932), .A2(net_931) );
CLKBUF_X2 inst_3070 ( .A(net_3027), .Z(net_3028) );
OAI21_X4 inst_85 ( .ZN(net_2046), .B1(net_2045), .A(net_2044), .B2(net_658) );
CLKBUF_X2 inst_2998 ( .A(net_2955), .Z(net_2956) );
CLKBUF_X2 inst_2916 ( .A(net_2873), .Z(net_2874) );
NAND2_X2 inst_1286 ( .A2(net_1858), .ZN(net_853), .A1(net_795) );
NOR2_X4 inst_266 ( .A2(net_2179), .ZN(net_1578), .A1(net_849) );
DFFR_X1 inst_2612 ( .Q(net_2772), .D(net_1845), .CK(net_2965), .RN(x2480) );
INV_X4 inst_2051 ( .ZN(net_1282), .A(net_1281) );
AOI22_X2 inst_2702 ( .A2(net_2759), .ZN(net_309), .B1(net_296), .A1(net_279), .B2(x1368) );
CLKBUF_X2 inst_2910 ( .A(net_2867), .Z(net_2868) );
NAND2_X2 inst_1198 ( .A1(net_1585), .A2(net_1533), .ZN(net_589) );
OAI21_X4 inst_77 ( .A(net_2557), .B2(net_2171), .B1(net_2014), .ZN(net_1739) );
OAI21_X2 inst_171 ( .ZN(net_2332), .B2(net_2331), .B1(net_2330), .A(net_2329) );
CLKBUF_X2 inst_3097 ( .A(net_2873), .Z(net_3055) );
NAND2_X2 inst_1362 ( .A1(net_2296), .A2(net_1559), .ZN(net_1152) );
CLKBUF_X2 inst_3238 ( .A(net_3195), .Z(net_3196) );
INV_X4 inst_1978 ( .A(net_2216), .ZN(net_805) );
OAI21_X2 inst_145 ( .ZN(net_1388), .B1(net_1387), .A(net_969), .B2(net_339) );
NOR2_X4 inst_290 ( .ZN(net_2087), .A2(net_2084), .A1(net_2083) );
NOR2_X2 inst_374 ( .A2(net_1843), .A1(net_1239), .ZN(net_788) );
NOR2_X4 inst_272 ( .A2(net_2360), .ZN(net_1718), .A1(net_1716) );
CLKBUF_X2 inst_3030 ( .A(net_2987), .Z(net_2988) );
CLKBUF_X2 inst_2854 ( .A(net_2811), .Z(net_2812) );
NAND4_X4 inst_502 ( .A2(net_1770), .ZN(net_1752), .A4(net_1751), .A1(net_1683), .A3(net_1053) );
INV_X4 inst_2112 ( .A(net_2567), .ZN(net_1915) );
OAI21_X4 inst_103 ( .ZN(net_2534), .A(net_2526), .B2(net_1360), .B1(net_505) );
CLKBUF_X2 inst_3036 ( .A(net_2993), .Z(net_2994) );
NAND2_X4 inst_814 ( .A1(net_2179), .ZN(net_1351), .A2(net_1312) );
INV_X2 inst_2230 ( .A(net_2433), .ZN(net_344) );
CLKBUF_X2 inst_3221 ( .A(net_3178), .Z(net_3179) );
NAND2_X2 inst_1458 ( .A1(net_2572), .ZN(net_1616), .A2(net_1615) );
INV_X2 inst_2275 ( .ZN(net_52), .A(x717) );
INV_X4 inst_1860 ( .A(net_1815), .ZN(net_485) );
INV_X8 inst_1810 ( .A(net_2647), .ZN(net_2129) );
INV_X8 inst_1806 ( .ZN(net_2062), .A(net_2052) );
NAND2_X4 inst_789 ( .ZN(net_1113), .A2(net_1112), .A1(net_1111) );
NAND2_X2 inst_1598 ( .ZN(net_2335), .A2(net_2334), .A1(net_2333) );
NOR2_X2 inst_357 ( .A2(net_2440), .A1(net_2357), .ZN(net_435) );
CLKBUF_X2 inst_2855 ( .A(x3333), .Z(net_2813) );
INV_X4 inst_1885 ( .A(net_1509), .ZN(net_363) );
NAND2_X2 inst_1437 ( .ZN(net_1444), .A1(net_1443), .A2(net_1142) );
INV_X4 inst_2058 ( .A(net_2288), .ZN(net_1352) );
NAND2_X4 inst_809 ( .A1(net_1658), .ZN(net_1311), .A2(net_1130) );
CLKBUF_X2 inst_3152 ( .A(net_2848), .Z(net_3110) );
NAND2_X4 inst_822 ( .ZN(net_1410), .A1(net_1409), .A2(net_1096) );
NAND2_X2 inst_1125 ( .A2(net_617), .A1(net_234), .ZN(net_213) );
DFFR_X1 inst_2562 ( .QN(net_2789), .Q(net_1479), .D(net_1328), .CK(net_3078), .RN(x2480) );
NAND2_X2 inst_1234 ( .A1(net_2489), .A2(net_1611), .ZN(net_657) );
NAND2_X4 inst_912 ( .ZN(net_1994), .A2(net_1905), .A1(net_1362) );
NAND3_X2 inst_609 ( .A2(net_1696), .ZN(net_1101), .A1(net_1099), .A3(net_918) );
INV_X2 inst_2398 ( .ZN(net_2513), .A(net_2512) );
DFFR_X1 inst_2595 ( .D(net_2770), .CK(net_3363), .RN(x2480), .Q(x258) );
NAND2_X4 inst_1022 ( .ZN(net_2631), .A1(net_2186), .A2(net_1906) );
DFFR_X2 inst_2533 ( .QN(net_2804), .D(net_85), .CK(net_3103), .RN(x2480) );
INV_X2 inst_2391 ( .ZN(net_2313), .A(net_2312) );
CLKBUF_X2 inst_3196 ( .A(net_3153), .Z(net_3154) );
DFFR_X2 inst_2496 ( .D(net_2459), .Q(net_1490), .CK(net_2962), .RN(x2480) );
INV_X2 inst_2371 ( .A(net_2031), .ZN(net_1818) );
NAND2_X4 inst_795 ( .A2(net_2179), .ZN(net_1192), .A1(net_849) );
INV_X2 inst_2239 ( .A(net_721), .ZN(net_327) );
OAI22_X2 inst_27 ( .B2(net_2286), .A2(net_2120), .A1(net_1548), .ZN(net_1239), .B1(net_571) );
CLKBUF_X2 inst_2939 ( .A(net_2896), .Z(net_2897) );
DFFR_X2 inst_2491 ( .Q(net_1499), .D(net_323), .CK(net_2866), .RN(x2480) );
NAND2_X2 inst_1639 ( .ZN(net_2571), .A1(net_2488), .A2(net_915) );
NOR2_X4 inst_322 ( .ZN(net_2564), .A1(net_2095), .A2(net_1725) );
NAND2_X2 inst_1223 ( .A1(net_1585), .A2(net_1490), .ZN(net_639) );
AOI21_X2 inst_2785 ( .B2(net_2250), .A(net_817), .ZN(net_466), .B1(net_402) );
NAND3_X2 inst_619 ( .A2(net_2590), .A1(net_1829), .ZN(net_1317), .A3(net_1316) );
NAND3_X2 inst_681 ( .ZN(net_2539), .A1(net_2528), .A2(net_1803), .A3(net_923) );
INV_X4 inst_2010 ( .A(net_2493), .ZN(net_1006) );
NAND2_X2 inst_1654 ( .ZN(net_2616), .A1(net_1850), .A2(net_957) );
CLKBUF_X2 inst_2915 ( .A(net_2872), .Z(net_2873) );
NAND2_X2 inst_1355 ( .ZN(net_1117), .A1(net_586), .A2(net_246) );
NAND3_X2 inst_639 ( .A3(net_2293), .ZN(net_1682), .A1(net_1333), .A2(net_992) );
NAND2_X4 inst_877 ( .A1(net_1878), .ZN(net_1796), .A2(net_178) );
CLKBUF_X2 inst_3296 ( .A(net_2848), .Z(net_3254) );
OAI21_X2 inst_155 ( .ZN(net_1763), .B1(net_156), .A(net_135), .B2(net_51) );
NAND2_X4 inst_871 ( .ZN(net_1765), .A2(net_1764), .A1(net_1762) );
INV_X2 inst_2315 ( .A(net_2055), .ZN(net_821) );
NAND2_X4 inst_962 ( .ZN(net_2289), .A2(net_2288), .A1(net_2287) );
NAND4_X2 inst_532 ( .A2(net_2562), .A3(net_2398), .A1(net_1916), .ZN(net_1729), .A4(net_809) );
OAI21_X4 inst_55 ( .B1(net_1585), .ZN(net_629), .A(net_132), .B2(net_41) );
CLKBUF_X2 inst_3164 ( .A(net_3051), .Z(net_3122) );
CLKBUF_X2 inst_2965 ( .A(net_2856), .Z(net_2923) );
INV_X2 inst_2382 ( .ZN(net_2031), .A(net_2030) );
INV_X2 inst_2280 ( .ZN(net_47), .A(x1611) );
INV_X4 inst_2167 ( .ZN(net_2441), .A(net_2440) );
INV_X4 inst_2008 ( .A(net_1364), .ZN(net_980) );
NAND2_X2 inst_1171 ( .ZN(net_564), .A1(net_86), .A2(x935) );
NAND3_X2 inst_641 ( .A2(net_1810), .ZN(net_1748), .A3(net_1221), .A1(net_1166) );
CLKBUF_X2 inst_2969 ( .A(net_2926), .Z(net_2927) );
NAND4_X4 inst_498 ( .A1(net_1187), .A3(net_1171), .A2(net_1157), .ZN(net_1017), .A4(net_879) );
CLKBUF_X2 inst_3314 ( .A(net_2861), .Z(net_3272) );
INV_X4 inst_1988 ( .ZN(net_845), .A(net_456) );
INV_X4 inst_2076 ( .ZN(net_1600), .A(net_1148) );
DFFR_X1 inst_2594 ( .D(net_2757), .CK(net_3146), .RN(x2480), .Q(x467) );
NAND2_X2 inst_1651 ( .ZN(net_2605), .A2(net_2604), .A1(net_1292) );
DFFR_X2 inst_2481 ( .Q(net_1516), .D(net_332), .CK(net_2880), .RN(x2480) );
INV_X4 inst_1912 ( .A(net_1514), .ZN(net_250) );
INV_X8 inst_1831 ( .ZN(net_2405), .A(net_2404) );
NAND2_X2 inst_1327 ( .A2(net_1641), .ZN(net_979), .A1(net_719) );
NAND2_X2 inst_1137 ( .A2(net_2320), .A1(net_617), .ZN(net_194) );
NOR2_X4 inst_323 ( .ZN(net_2568), .A2(net_347), .A1(net_341) );
NAND2_X2 inst_1162 ( .A2(net_1505), .ZN(net_118), .A1(net_117) );
NAND2_X2 inst_1389 ( .ZN(net_1273), .A1(net_498), .A2(net_492) );
NOR2_X2 inst_350 ( .A2(net_2165), .A1(net_1790), .ZN(net_419) );
CLKBUF_X2 inst_2973 ( .A(net_2930), .Z(net_2931) );
INV_X2 inst_2395 ( .ZN(net_2444), .A(net_2440) );
NOR2_X4 inst_231 ( .ZN(net_997), .A1(net_273), .A2(net_256) );
CLKBUF_X2 inst_3065 ( .A(net_3022), .Z(net_3023) );
NAND2_X2 inst_1119 ( .A1(net_1191), .A2(net_234), .ZN(net_223) );
NAND2_X2 inst_1494 ( .ZN(net_1757), .A1(net_116), .A2(net_100) );
NAND2_X2 inst_1433 ( .A1(net_2691), .ZN(net_1404), .A2(net_744) );
NAND2_X4 inst_793 ( .ZN(net_1191), .A2(net_1190), .A1(net_587) );
NAND2_X4 inst_715 ( .A1(net_1410), .A2(net_221), .ZN(net_175) );
CLKBUF_X2 inst_3309 ( .A(net_3266), .Z(net_3267) );
INV_X4 inst_1894 ( .A(net_2398), .ZN(net_346) );
NAND2_X2 inst_1255 ( .A2(net_2111), .A1(net_1194), .ZN(net_731) );
CLKBUF_X2 inst_3449 ( .A(net_3406), .Z(net_3407) );
INV_X2 inst_2317 ( .A(net_1167), .ZN(net_872) );
INV_X4 inst_1999 ( .ZN(net_929), .A(net_928) );
NAND2_X2 inst_1682 ( .ZN(net_2735), .A2(net_2106), .A1(net_2105) );
AOI22_X2 inst_2733 ( .A2(net_2751), .ZN(net_1969), .B1(net_296), .A1(net_283), .B2(x1405) );
NAND2_X2 inst_1481 ( .A1(net_2360), .ZN(net_1724), .A2(net_1722) );
NAND2_X2 inst_1340 ( .A2(net_1236), .ZN(net_1046), .A1(net_570) );
INV_X8 inst_1791 ( .A(net_1824), .ZN(net_1822) );
NAND2_X2 inst_1452 ( .A2(net_2598), .ZN(net_1590), .A1(net_224) );
CLKBUF_X2 inst_3420 ( .A(net_3377), .Z(net_3378) );
NOR2_X2 inst_475 ( .ZN(net_2448), .A1(net_2447), .A2(net_1966) );
CLKBUF_X2 inst_3139 ( .A(net_3096), .Z(net_3097) );
AOI22_X2 inst_2701 ( .A2(net_2760), .ZN(net_310), .A1(net_279), .B1(net_278), .B2(x1517) );
OAI22_X2 inst_31 ( .B2(net_2786), .ZN(net_1978), .B1(net_633), .A1(net_143), .A2(net_45) );
NAND4_X2 inst_528 ( .ZN(net_1552), .A1(net_1551), .A2(net_903), .A3(net_702), .A4(net_512) );
DFFR_X1 inst_2558 ( .QN(net_2800), .Q(net_1522), .D(net_1019), .CK(net_3100), .RN(x2480) );
NAND2_X4 inst_903 ( .ZN(net_1960), .A2(net_1959), .A1(net_1957) );
CLKBUF_X2 inst_3165 ( .A(net_3036), .Z(net_3123) );
NAND2_X1 inst_1725 ( .A1(net_2129), .A2(net_1918), .ZN(net_1816) );
CLKBUF_X2 inst_3217 ( .A(net_3174), .Z(net_3175) );
NAND2_X2 inst_1396 ( .A1(net_2358), .A2(net_1546), .ZN(net_1296) );
NOR2_X2 inst_352 ( .A2(net_2153), .ZN(net_381), .A1(net_359) );
NAND3_X4 inst_575 ( .ZN(net_2201), .A1(net_2200), .A2(net_271), .A3(net_208) );
NAND2_X4 inst_846 ( .ZN(net_1623), .A1(net_1044), .A2(net_364) );
NOR2_X4 inst_286 ( .A2(net_2157), .ZN(net_2027), .A1(net_2026) );
INV_X8 inst_1734 ( .ZN(net_385), .A(net_367) );
NAND3_X2 inst_627 ( .ZN(net_1545), .A1(net_1544), .A3(net_979), .A2(net_978) );
CLKBUF_X2 inst_3352 ( .A(net_3309), .Z(net_3310) );
NOR2_X2 inst_344 ( .A2(net_2137), .A1(net_435), .ZN(net_423) );
INV_X8 inst_1833 ( .A(net_2611), .ZN(net_2426) );
CLKBUF_X2 inst_3044 ( .A(net_3001), .Z(net_3002) );
INV_X4 inst_2122 ( .ZN(net_1988), .A(net_1987) );
CLKBUF_X2 inst_3003 ( .A(net_2960), .Z(net_2961) );
CLKBUF_X2 inst_3464 ( .A(net_3057), .Z(net_3422) );
INV_X4 inst_2185 ( .ZN(net_2622), .A(net_2621) );
NAND3_X2 inst_623 ( .A2(net_2178), .ZN(net_1914), .A3(net_933), .A1(net_655) );
NAND2_X2 inst_1072 ( .A2(net_2061), .A1(net_707), .ZN(net_477) );
NAND2_X2 inst_1044 ( .A1(net_2332), .A2(net_2142), .ZN(net_561) );
CLKBUF_X2 inst_3354 ( .A(net_3311), .Z(net_3312) );
INV_X4 inst_1993 ( .A(net_936), .ZN(net_864) );
NAND2_X2 inst_1621 ( .ZN(net_2468), .A2(net_2464), .A1(net_1428) );
NAND2_X2 inst_1338 ( .A2(net_2414), .ZN(net_1022), .A1(net_764) );
INV_X16 inst_2430 ( .ZN(net_2259), .A(net_86) );
INV_X2 inst_2370 ( .ZN(net_1783), .A(net_1782) );
CLKBUF_X2 inst_3080 ( .A(net_3037), .Z(net_3038) );
INV_X16 inst_2434 ( .ZN(net_2360), .A(net_2359) );
CLKBUF_X2 inst_3226 ( .A(net_2946), .Z(net_3184) );
NAND2_X2 inst_1107 ( .A2(net_660), .ZN(net_268), .A1(net_215) );
AOI21_X2 inst_2811 ( .ZN(net_1872), .B1(net_1870), .A(net_1181), .B2(net_822) );
INV_X4 inst_2028 ( .ZN(net_1127), .A(net_1126) );
NAND2_X2 inst_1377 ( .A1(net_2655), .ZN(net_1210), .A2(net_736) );
CLKBUF_X2 inst_3014 ( .A(net_2971), .Z(net_2972) );
CLKBUF_X2 inst_3125 ( .A(net_3082), .Z(net_3083) );
INV_X2 inst_2201 ( .A(net_993), .ZN(net_516) );
OAI21_X2 inst_137 ( .B1(net_2390), .B2(net_1799), .ZN(net_1144), .A(net_490) );
NOR2_X2 inst_425 ( .A1(net_2726), .A2(net_2136), .ZN(net_1387) );
DFFR_X1 inst_2567 ( .D(net_2780), .CK(net_2859), .RN(x2480), .Q(x363) );
CLKBUF_X2 inst_3206 ( .A(net_2957), .Z(net_3164) );
AOI21_X4 inst_2776 ( .A(net_2397), .ZN(net_2090), .B1(net_1063), .B2(net_681) );
NAND2_X2 inst_1532 ( .ZN(net_1986), .A1(net_1985), .A2(x1851) );
NAND2_X4 inst_722 ( .A2(net_1213), .A1(net_1212), .ZN(net_203) );
NOR2_X4 inst_227 ( .A1(net_1101), .A2(net_1066), .ZN(net_913) );
NAND2_X4 inst_760 ( .A1(net_2731), .A2(net_2099), .ZN(net_841) );
INV_X4 inst_2136 ( .ZN(net_2145), .A(net_2143) );
NAND2_X4 inst_746 ( .A1(net_2739), .ZN(net_717), .A2(net_716) );
CLKBUF_X2 inst_2891 ( .A(net_2848), .Z(net_2849) );
AOI22_X2 inst_2718 ( .B1(net_883), .ZN(net_855), .B2(net_854), .A2(net_852), .A1(net_851) );
DFFR_X1 inst_2572 ( .D(net_2764), .CK(net_2903), .RN(x2480), .Q(x397) );
OAI21_X4 inst_58 ( .B1(net_1585), .ZN(net_647), .A(net_646), .B2(net_48) );
NAND2_X1 inst_1696 ( .ZN(net_231), .A2(net_217), .A1(net_187) );
INV_X2 inst_2267 ( .ZN(net_60), .A(x1312) );
CLKBUF_X2 inst_3010 ( .A(net_2967), .Z(net_2968) );
CLKBUF_X2 inst_3365 ( .A(net_3322), .Z(net_3323) );
NAND2_X2 inst_1469 ( .A2(net_2293), .ZN(net_1680), .A1(net_902) );
CLKBUF_X2 inst_3254 ( .A(net_3211), .Z(net_3212) );
NAND2_X4 inst_983 ( .ZN(net_2390), .A1(net_1646), .A2(net_361) );
CLKBUF_X2 inst_3133 ( .A(net_3090), .Z(net_3091) );
INV_X4 inst_1897 ( .ZN(net_394), .A(net_342) );
CLKBUF_X2 inst_3159 ( .A(net_3116), .Z(net_3117) );
NAND2_X1 inst_1687 ( .A1(net_527), .A2(net_472), .ZN(net_462) );
NAND2_X2 inst_1577 ( .ZN(net_2194), .A1(net_2193), .A2(net_2107) );
DFFR_X1 inst_2588 ( .Q(net_2760), .D(net_1514), .CK(net_3262), .RN(x2480) );
DFFR_X1 inst_2551 ( .QN(net_2793), .Q(net_1487), .D(net_897), .CK(net_3279), .RN(x2480) );
INV_X4 inst_1970 ( .A(net_813), .ZN(net_764) );
NAND2_X2 inst_1110 ( .A2(net_1734), .ZN(net_258), .A1(net_188) );
NAND3_X4 inst_581 ( .ZN(net_2497), .A2(net_2496), .A3(net_2495), .A1(net_2494) );
OAI22_X2 inst_28 ( .ZN(net_1313), .A1(net_1078), .A2(net_817), .B2(net_527), .B1(net_467) );
INV_X16 inst_2424 ( .ZN(net_2111), .A(net_2110) );
CLKBUF_X2 inst_2873 ( .A(net_2813), .Z(net_2831) );
NAND2_X2 inst_1569 ( .ZN(net_2155), .A1(net_1329), .A2(net_607) );
INV_X16 inst_2442 ( .ZN(net_2561), .A(net_2560) );
CLKBUF_X2 inst_3144 ( .A(net_3101), .Z(net_3102) );
DFFR_X1 inst_2633 ( .D(net_75), .CK(net_3393), .RN(x2480), .Q(x279) );
INV_X8 inst_1772 ( .A(net_2433), .ZN(net_1167) );
NAND3_X2 inst_592 ( .A1(net_737), .ZN(net_272), .A3(net_230), .A2(net_197) );
CLKBUF_X2 inst_3411 ( .A(net_3368), .Z(net_3369) );
INV_X4 inst_2066 ( .ZN(net_1461), .A(net_1460) );
NAND2_X4 inst_993 ( .ZN(net_2460), .A1(net_2459), .A2(net_152) );
INV_X4 inst_2143 ( .ZN(net_2222), .A(net_2220) );
DFFR_X2 inst_2524 ( .D(net_1957), .Q(net_1496), .CK(net_3109), .RN(x2480) );
NAND2_X2 inst_1446 ( .ZN(net_1557), .A2(net_1556), .A1(net_1555) );
NAND2_X2 inst_1291 ( .A2(net_2533), .ZN(net_874), .A1(net_829) );
INV_X16 inst_2421 ( .ZN(net_2061), .A(net_1715) );
NOR2_X2 inst_390 ( .A2(net_1167), .ZN(net_938), .A1(net_382) );
INV_X8 inst_1742 ( .A(net_1073), .ZN(net_340) );
INV_X4 inst_2130 ( .ZN(net_2059), .A(net_2058) );
NAND2_X2 inst_1062 ( .A1(net_2406), .A2(net_1035), .ZN(net_506) );
NOR2_X2 inst_359 ( .A1(net_2408), .A2(net_1429), .ZN(net_357) );
NAND2_X2 inst_1055 ( .A1(net_1995), .A2(net_718), .ZN(net_531) );
CLKBUF_X2 inst_3289 ( .A(net_2997), .Z(net_3247) );
CLKBUF_X2 inst_2875 ( .A(net_2832), .Z(net_2833) );
DFFR_X1 inst_2663 ( .D(net_1471), .CK(net_3359), .RN(x2480), .Q(x253) );
INV_X4 inst_2100 ( .ZN(net_1795), .A(net_1313) );
INV_X2 inst_2284 ( .ZN(net_43), .A(x1800) );
INV_X4 inst_1962 ( .A(net_2138), .ZN(net_708) );
NAND3_X2 inst_630 ( .A2(net_2567), .A1(net_2393), .A3(net_1725), .ZN(net_1572) );
CLKBUF_X2 inst_3175 ( .A(net_2849), .Z(net_3133) );
INV_X2 inst_2302 ( .ZN(net_599), .A(x1007) );
NOR2_X2 inst_401 ( .A1(net_2215), .A2(net_1678), .ZN(net_1042) );
NAND2_X2 inst_1273 ( .ZN(net_784), .A2(net_227), .A1(net_187) );
CLKBUF_X2 inst_3389 ( .A(net_3346), .Z(net_3347) );
NAND2_X4 inst_923 ( .ZN(net_2052), .A1(net_337), .A2(net_336) );
NAND4_X2 inst_512 ( .A2(net_1763), .ZN(net_751), .A1(net_311), .A3(net_269), .A4(net_253) );
CLKBUF_X2 inst_3210 ( .A(net_3167), .Z(net_3168) );
INV_X1 inst_2447 ( .A(net_1176), .ZN(net_652) );
NAND2_X2 inst_1301 ( .ZN(net_900), .A1(net_521), .A2(net_482) );
NAND2_X4 inst_782 ( .ZN(net_1076), .A1(net_1075), .A2(net_640) );
INV_X4 inst_2151 ( .ZN(net_2326), .A(net_2325) );
AND2_X4 inst_2830 ( .ZN(net_1890), .A1(net_1425), .A2(net_1423) );
NAND3_X2 inst_647 ( .A3(net_2738), .ZN(net_1923), .A1(net_1907), .A2(net_1362) );
CLKBUF_X2 inst_3054 ( .A(net_3011), .Z(net_3012) );
DFFR_X1 inst_2642 ( .D(net_74), .CK(net_3242), .RN(x2480), .Q(x121) );
CLKBUF_X2 inst_2869 ( .A(net_2819), .Z(net_2827) );
OR2_X4 inst_6 ( .ZN(net_2455), .A2(net_2454), .A1(net_2453) );
NOR3_X4 inst_194 ( .A2(net_1335), .A3(net_714), .ZN(net_487), .A1(net_427) );
DFFR_X2 inst_2486 ( .Q(net_1528), .D(net_320), .CK(net_2875), .RN(x2480) );
CLKBUF_X2 inst_3453 ( .A(net_3174), .Z(net_3411) );
CLKBUF_X2 inst_2985 ( .A(net_2942), .Z(net_2943) );
INV_X16 inst_2410 ( .A(net_658), .ZN(net_586) );
NAND2_X4 inst_833 ( .A1(net_1767), .ZN(net_1546), .A2(net_367) );
OAI21_X2 inst_123 ( .B1(net_1690), .ZN(net_814), .B2(net_255), .A(net_213) );
NAND2_X4 inst_930 ( .ZN(net_2104), .A1(net_722), .A2(net_579) );
DFFR_X1 inst_2536 ( .QN(net_2782), .Q(net_1501), .D(net_1398), .CK(net_3253), .RN(x2480) );
INV_X4 inst_2043 ( .ZN(net_1232), .A(net_1231) );
NAND2_X4 inst_960 ( .ZN(net_2277), .A1(net_2276), .A2(net_1757) );
OAI21_X2 inst_118 ( .B1(net_1335), .A(net_849), .ZN(net_611), .B2(net_407) );
INV_X4 inst_2160 ( .ZN(net_2393), .A(net_2392) );
INV_X16 inst_2411 ( .A(net_1585), .ZN(net_635) );
NAND2_X4 inst_935 ( .ZN(net_2134), .A2(net_2133), .A1(net_2131) );
NOR2_X2 inst_442 ( .A1(net_2429), .A2(net_1822), .ZN(net_1679) );
DFFR_X2 inst_2507 ( .D(net_2088), .Q(net_1481), .CK(net_3210), .RN(x2480) );
INV_X2 inst_2245 ( .A(net_622), .ZN(net_170) );
OAI221_X2 inst_38 ( .C2(net_1690), .ZN(net_324), .B2(net_319), .A(net_305), .B1(net_181), .C1(net_145) );
DFFR_X1 inst_2601 ( .Q(net_2751), .D(net_2106), .CK(net_3347), .RN(x2480) );
INV_X4 inst_2037 ( .ZN(net_1185), .A(net_1184) );
NOR2_X2 inst_381 ( .A2(net_2737), .A1(net_2453), .ZN(net_875) );
INV_X2 inst_2298 ( .ZN(net_30), .A(x554) );
INV_X4 inst_1925 ( .A(net_182), .ZN(net_160) );
NAND2_X4 inst_883 ( .ZN(net_1837), .A1(net_1585), .A2(net_1489) );
OAI221_X2 inst_40 ( .C2(net_857), .ZN(net_322), .C1(net_321), .B2(net_319), .A(net_304), .B1(net_193) );
NAND2_X2 inst_1249 ( .A2(net_1907), .ZN(net_719), .A1(net_716) );
OAI21_X2 inst_167 ( .A(net_2546), .ZN(net_2298), .B2(net_2297), .B1(net_2293) );
CLKBUF_X2 inst_2944 ( .A(net_2901), .Z(net_2902) );
NAND2_X2 inst_1320 ( .A2(net_2133), .ZN(net_964), .A1(net_209) );
NAND2_X4 inst_1026 ( .ZN(net_2655), .A1(net_624), .A2(net_92) );
NAND2_X4 inst_756 ( .ZN(net_794), .A2(net_493), .A1(net_401) );
NAND2_X2 inst_1251 ( .ZN(net_723), .A1(net_721), .A2(net_209) );
CLKBUF_X2 inst_3376 ( .A(net_3333), .Z(net_3334) );
NAND2_X2 inst_1416 ( .A1(net_2279), .ZN(net_1350), .A2(net_314) );
OAI21_X4 inst_95 ( .ZN(net_2262), .B2(net_2261), .A(net_2260), .B1(net_2259) );
DFFR_X2 inst_2475 ( .D(net_1762), .Q(net_1519), .CK(net_3117), .RN(x2480) );
NAND2_X2 inst_1318 ( .ZN(net_962), .A2(net_961), .A1(net_778) );
CLKBUF_X2 inst_2921 ( .A(net_2878), .Z(net_2879) );
NOR2_X2 inst_439 ( .ZN(net_1627), .A1(net_1626), .A2(net_277) );
CLKBUF_X2 inst_2862 ( .A(net_2819), .Z(net_2820) );
NAND2_X2 inst_1188 ( .A2(net_2239), .ZN(net_2048), .A1(net_616) );
NAND2_X2 inst_1165 ( .A1(net_115), .ZN(net_111), .A2(net_72) );
NOR2_X4 inst_331 ( .ZN(net_2685), .A1(net_1710), .A2(net_261) );
DFFR_X1 inst_2644 ( .D(net_1487), .CK(net_3390), .RN(x2480), .Q(x266) );
NAND2_X2 inst_1070 ( .A1(net_1085), .A2(net_609), .ZN(net_480) );
DFFR_X1 inst_2626 ( .Q(net_2768), .D(net_179), .CK(net_3026), .RN(x2480) );
INV_X1 inst_2454 ( .A(net_243), .ZN(net_145) );
INV_X4 inst_2172 ( .ZN(net_2494), .A(net_1755) );
INV_X2 inst_2353 ( .ZN(net_1586), .A(net_1585) );
NAND3_X2 inst_667 ( .A3(net_2338), .ZN(net_2220), .A1(net_1601), .A2(net_504) );
AOI21_X4 inst_2762 ( .B2(net_1215), .B1(net_1214), .A(net_937), .ZN(net_839) );
NAND2_X4 inst_992 ( .ZN(net_2453), .A1(net_2109), .A2(net_1913) );
NOR2_X2 inst_488 ( .ZN(net_2729), .A2(net_2647), .A1(net_2562) );
CLKBUF_X2 inst_2896 ( .A(net_2853), .Z(net_2854) );
NOR2_X2 inst_387 ( .ZN(net_923), .A1(net_922), .A2(net_921) );
NAND2_X4 inst_997 ( .A1(net_2489), .ZN(net_2469), .A2(net_1738) );
NAND2_X4 inst_857 ( .A1(net_2284), .ZN(net_1684), .A2(net_350) );
NOR2_X4 inst_254 ( .A2(net_1905), .ZN(net_1361), .A1(net_1359) );
NAND3_X2 inst_654 ( .ZN(net_1967), .A2(net_1795), .A1(net_1794), .A3(net_1058) );
AOI22_X4 inst_2691 ( .B1(net_2309), .A2(net_1859), .ZN(net_1049), .A1(net_1048), .B2(net_854) );
NAND2_X2 inst_1673 ( .ZN(net_2704), .A2(net_955), .A1(net_476) );
NAND2_X2 inst_1511 ( .ZN(net_1875), .A1(net_1874), .A2(net_744) );
INV_X4 inst_2129 ( .ZN(net_2045), .A(net_266) );
NAND2_X2 inst_1412 ( .A1(net_2605), .ZN(net_1342), .A2(net_309) );
NOR2_X2 inst_365 ( .A2(net_2165), .A1(net_2061), .ZN(net_608) );
NAND2_X1 inst_1708 ( .ZN(net_706), .A2(net_705), .A1(net_704) );
NAND2_X2 inst_1181 ( .ZN(net_2733), .A1(net_86), .A2(x692) );
OAI21_X4 inst_67 ( .B1(net_2592), .ZN(net_1233), .A(net_741), .B2(net_233) );
CLKBUF_X2 inst_3203 ( .A(net_2866), .Z(net_3161) );
NAND2_X4 inst_954 ( .ZN(net_2235), .A1(net_2234), .A2(net_929) );
NAND2_X2 inst_1153 ( .A2(net_1540), .ZN(net_131), .A1(net_130) );
NAND2_X2 inst_1504 ( .ZN(net_1841), .A1(net_1840), .A2(net_1355) );
DFFR_X2 inst_2476 ( .Q(net_1507), .D(net_1118), .CK(net_3255), .RN(x2480) );
NOR2_X2 inst_391 ( .A2(net_2803), .ZN(net_941), .A1(net_81) );
CLKBUF_X2 inst_3403 ( .A(net_3290), .Z(net_3361) );
NAND3_X2 inst_661 ( .ZN(net_2103), .A3(net_734), .A2(net_567), .A1(net_566) );
INV_X8 inst_1823 ( .ZN(net_2325), .A(net_2320) );
NAND2_X2 inst_1548 ( .ZN(net_2077), .A1(net_2068), .A2(net_1611) );
INV_X4 inst_2073 ( .ZN(net_1581), .A(net_1579) );
NAND2_X2 inst_1310 ( .A2(net_2603), .A1(net_1167), .ZN(net_936) );
NOR3_X2 inst_202 ( .A3(net_2726), .A1(net_2444), .A2(net_2288), .ZN(net_1426) );
INV_X2 inst_2212 ( .A(net_2577), .ZN(net_412) );
CLKBUF_X2 inst_3280 ( .A(net_3237), .Z(net_3238) );
NAND2_X2 inst_1401 ( .A1(net_1658), .ZN(net_1312), .A2(net_1130) );
AOI22_X2 inst_2738 ( .ZN(net_2316), .B2(net_2239), .A2(net_647), .A1(net_586), .B1(net_216) );
NAND3_X2 inst_634 ( .ZN(net_1633), .A1(net_1266), .A3(net_770), .A2(net_543) );
NOR2_X2 inst_419 ( .ZN(net_1343), .A1(net_1273), .A2(net_896) );
CLKBUF_X2 inst_3122 ( .A(net_3079), .Z(net_3080) );
AND4_X4 inst_2823 ( .A2(net_2495), .ZN(net_1759), .A4(net_1758), .A3(net_1757), .A1(net_1756) );
INV_X4 inst_2030 ( .ZN(net_1146), .A(net_1145) );
NAND2_X2 inst_1069 ( .A1(net_1332), .ZN(net_482), .A2(net_368) );
OAI21_X2 inst_136 ( .B2(net_1285), .A(net_1218), .ZN(net_1135), .B1(net_1034) );
OAI22_X2 inst_30 ( .A2(net_2285), .ZN(net_1843), .A1(net_1437), .B1(net_1320), .B2(net_685) );
NAND3_X2 inst_610 ( .A2(net_2129), .A3(net_1915), .ZN(net_1138), .A1(net_437) );
NAND2_X4 inst_1036 ( .ZN(net_2716), .A1(net_1879), .A2(net_1106) );
NOR2_X4 inst_233 ( .A1(net_1144), .ZN(net_1036), .A2(net_891) );
NAND2_X2 inst_1526 ( .ZN(net_1958), .A1(net_120), .A2(net_106) );
NAND2_X2 inst_1477 ( .ZN(net_1708), .A2(net_1689), .A1(net_927) );
DFFR_X1 inst_2547 ( .D(net_2451), .Q(net_71), .CK(net_2924), .RN(x2480) );
OAI22_X2 inst_34 ( .B1(net_2493), .ZN(net_2474), .A1(net_2469), .B2(net_2070), .A2(net_1611) );
INV_X8 inst_1799 ( .ZN(net_1913), .A(net_1912) );
OR2_X2 inst_12 ( .A2(net_2800), .ZN(net_1330), .A1(net_634) );
NAND2_X2 inst_1047 ( .A2(net_750), .ZN(net_555), .A1(net_531) );
NAND4_X2 inst_529 ( .ZN(net_1592), .A2(net_1591), .A3(net_689), .A1(net_267), .A4(net_182) );
NAND2_X2 inst_1528 ( .A1(net_2602), .ZN(net_1971), .A2(net_936) );
OAI21_X4 inst_60 ( .B2(net_2406), .A(net_2339), .ZN(net_865), .B1(net_533) );
CLKBUF_X2 inst_3458 ( .A(net_3415), .Z(net_3416) );
NAND2_X2 inst_1424 ( .A2(net_1689), .A1(net_1577), .ZN(net_1380) );
INV_X4 inst_1858 ( .A(net_583), .ZN(net_469) );
INV_X8 inst_1786 ( .A(net_2351), .ZN(net_1720) );
NAND2_X2 inst_1313 ( .A1(net_1904), .A2(net_1510), .ZN(net_949) );
INV_X2 inst_2376 ( .ZN(net_1856), .A(net_1855) );
NAND2_X2 inst_1425 ( .A2(net_2237), .A1(net_1577), .ZN(net_1381) );
NAND2_X2 inst_1334 ( .A2(net_2312), .A1(net_1903), .ZN(net_1002) );
NAND3_X2 inst_675 ( .ZN(net_2400), .A3(net_2399), .A2(net_2397), .A1(net_2393) );
NOR2_X1 inst_496 ( .ZN(net_2742), .A2(net_1359), .A1(net_717) );
NAND2_X4 inst_860 ( .ZN(net_1694), .A2(net_1693), .A1(net_1692) );
CLKBUF_X2 inst_2886 ( .A(net_2840), .Z(net_2844) );
NAND4_X1 inst_563 ( .A3(net_2543), .ZN(net_2529), .A1(net_2528), .A2(net_1803), .A4(net_920) );
AOI22_X2 inst_2705 ( .A2(net_2764), .ZN(net_307), .A1(net_295), .B1(net_126), .B2(x1993) );
INV_X2 inst_2307 ( .ZN(net_773), .A(net_222) );
INV_X4 inst_2198 ( .ZN(net_2746), .A(net_2745) );
NAND2_X4 inst_943 ( .A1(net_2282), .ZN(net_2175), .A2(net_1350) );
NOR2_X4 inst_258 ( .A2(net_1644), .ZN(net_1420), .A1(net_657) );
DFFR_X1 inst_2611 ( .Q(net_2761), .D(net_1763), .CK(net_3345), .RN(x2480) );
AOI21_X4 inst_2773 ( .ZN(net_1773), .A(net_1386), .B2(net_836), .B1(net_544) );
INV_X4 inst_2081 ( .ZN(net_1646), .A(net_1644) );
CLKBUF_X2 inst_3261 ( .A(net_3218), .Z(net_3219) );
DFFR_X1 inst_2620 ( .Q(net_2755), .D(net_1978), .CK(net_3091), .RN(x2480) );
INV_X2 inst_2405 ( .ZN(net_2659), .A(net_1854) );
AOI21_X2 inst_2782 ( .B2(net_2022), .A(net_853), .ZN(net_548), .B1(net_487) );
CLKBUF_X2 inst_2994 ( .A(net_2854), .Z(net_2952) );
INV_X4 inst_1964 ( .ZN(net_718), .A(net_716) );
CLKBUF_X2 inst_3023 ( .A(net_2980), .Z(net_2981) );
INV_X8 inst_1765 ( .A(net_1311), .ZN(net_849) );
NAND2_X2 inst_1633 ( .ZN(net_2535), .A2(net_2525), .A1(net_2512) );
NAND2_X2 inst_1262 ( .A1(net_2133), .A2(net_1469), .ZN(net_741) );
NAND2_X2 inst_1243 ( .A2(net_2320), .ZN(net_687), .A1(net_212) );
NOR2_X4 inst_265 ( .A2(net_2027), .ZN(net_1561), .A1(net_1560) );
CLKBUF_X2 inst_3076 ( .A(net_3033), .Z(net_3034) );
INV_X4 inst_2055 ( .ZN(net_1302), .A(net_1299) );
INV_X4 inst_2005 ( .ZN(net_961), .A(net_959) );
NAND2_X2 inst_1211 ( .A1(net_1585), .A2(net_1464), .ZN(net_623) );
NOR2_X2 inst_482 ( .ZN(net_2572), .A2(net_2071), .A1(net_1070) );
NAND2_X2 inst_1192 ( .A1(net_2386), .A2(net_1448), .ZN(net_578) );
NAND3_X2 inst_682 ( .ZN(net_2546), .A1(net_2545), .A2(net_1927), .A3(net_1820) );
NAND2_X4 inst_736 ( .A1(net_1585), .A2(net_1526), .ZN(net_591) );
NAND4_X2 inst_544 ( .A3(net_2583), .ZN(net_2064), .A2(net_2063), .A4(net_2062), .A1(net_2061) );
NOR2_X4 inst_238 ( .A2(net_2582), .ZN(net_1108), .A1(net_1107) );
CLKBUF_X2 inst_3276 ( .A(net_3089), .Z(net_3234) );
NAND2_X2 inst_1093 ( .A2(net_2178), .A1(net_1335), .ZN(net_376) );
NAND4_X2 inst_539 ( .A2(net_1958), .A1(net_1956), .ZN(net_1881), .A4(net_726), .A3(net_184) );
INV_X2 inst_2222 ( .A(net_817), .ZN(net_365) );
CLKBUF_X2 inst_3333 ( .A(net_2843), .Z(net_3291) );
CLKBUF_X2 inst_3262 ( .A(net_3219), .Z(net_3220) );
NAND2_X4 inst_895 ( .ZN(net_1933), .A2(net_1932), .A1(net_1931) );
OAI21_X2 inst_178 ( .ZN(net_2638), .B2(net_2637), .B1(net_2634), .A(net_1173) );
CLKBUF_X2 inst_3109 ( .A(net_3066), .Z(net_3067) );
CLKBUF_X2 inst_3271 ( .A(net_3228), .Z(net_3229) );
NAND2_X2 inst_1430 ( .ZN(net_1389), .A2(net_948), .A1(net_947) );
NAND2_X4 inst_734 ( .A2(net_2267), .A1(net_769), .ZN(net_583) );
INV_X8 inst_1755 ( .ZN(net_598), .A(net_98) );
CLKBUF_X2 inst_3257 ( .A(net_3214), .Z(net_3215) );
INV_X2 inst_2240 ( .A(net_229), .ZN(net_220) );
NAND2_X2 inst_1282 ( .A2(net_2067), .A1(net_1610), .ZN(net_835) );
NAND2_X2 inst_1077 ( .A1(net_1163), .ZN(net_501), .A2(net_363) );
NAND2_X2 inst_1210 ( .A1(net_1585), .A2(net_1499), .ZN(net_620) );
INV_X2 inst_2341 ( .ZN(net_1326), .A(net_297) );
NAND2_X2 inst_1148 ( .A2(net_1564), .A1(net_180), .ZN(net_167) );
AOI222_X1 inst_2757 ( .A2(net_1877), .C2(net_1818), .C1(net_736), .ZN(net_735), .B1(net_721), .B2(net_220), .A1(net_158) );
INV_X16 inst_2437 ( .ZN(net_2396), .A(net_2395) );
INV_X4 inst_1932 ( .A(net_180), .ZN(net_159) );
NOR2_X4 inst_222 ( .ZN(net_796), .A2(net_795), .A1(net_794) );
NAND2_X4 inst_806 ( .A2(net_2404), .A1(net_1964), .ZN(net_1286) );
INV_X4 inst_1981 ( .ZN(net_817), .A(net_816) );
NAND2_X4 inst_763 ( .ZN(net_909), .A2(net_736), .A1(net_173) );
INV_X2 inst_2330 ( .ZN(net_1067), .A(net_1066) );
NOR2_X1 inst_491 ( .A2(net_1021), .ZN(net_800), .A1(net_385) );
NAND2_X2 inst_1302 ( .A1(net_1717), .ZN(net_902), .A2(net_805) );
NAND2_X2 inst_1280 ( .A2(net_1164), .A1(net_981), .ZN(net_829) );
NAND2_X2 inst_1052 ( .ZN(net_536), .A1(net_514), .A2(net_478) );
NAND2_X2 inst_1648 ( .ZN(net_2599), .A2(net_2597), .A1(net_187) );
NAND2_X2 inst_1079 ( .A2(net_986), .ZN(net_459), .A1(net_400) );
NAND2_X4 inst_842 ( .ZN(net_1602), .A1(net_626), .A2(net_96) );
NAND4_X2 inst_537 ( .ZN(net_1849), .A1(net_1848), .A3(net_1772), .A2(net_1771), .A4(net_831) );
INV_X4 inst_2068 ( .A(net_1680), .ZN(net_1551) );
INV_X1 inst_2472 ( .ZN(net_2502), .A(net_2501) );
NAND2_X4 inst_826 ( .A2(net_2137), .ZN(net_1437), .A1(net_961) );
CLKBUF_X2 inst_3086 ( .A(net_3043), .Z(net_3044) );
AOI21_X2 inst_2791 ( .B1(net_1859), .B2(net_846), .ZN(net_770), .A(net_466) );
DFFR_X1 inst_2606 ( .D(net_2766), .CK(net_3172), .RN(x2480), .Q(x31) );
NAND4_X2 inst_551 ( .ZN(net_2479), .A2(net_2476), .A1(net_1627), .A3(net_1094), .A4(net_552) );
DFFR_X2 inst_2523 ( .D(net_2201), .Q(net_1478), .CK(net_3285), .RN(x2480) );
INV_X4 inst_2101 ( .A(net_1965), .ZN(net_1797) );
NOR2_X2 inst_353 ( .A1(net_1567), .A2(net_1429), .ZN(net_377) );
NAND4_X4 inst_506 ( .ZN(net_2275), .A4(net_1210), .A1(net_1209), .A2(net_1091), .A3(net_195) );
OAI21_X2 inst_159 ( .B2(net_2789), .ZN(net_1987), .A(net_1986), .B1(net_225) );
NAND2_X4 inst_872 ( .ZN(net_1770), .A2(net_1769), .A1(net_1766) );
INV_X4 inst_1940 ( .A(net_1585), .ZN(net_169) );
CLKBUF_X2 inst_3322 ( .A(net_2829), .Z(net_3280) );
INV_X16 inst_2409 ( .A(net_1585), .ZN(net_86) );
OAI21_X2 inst_134 ( .A(net_2165), .B1(net_2156), .B2(net_2065), .ZN(net_1109) );
CLKBUF_X2 inst_3425 ( .A(net_3382), .Z(net_3383) );
NAND2_X2 inst_1323 ( .A1(net_1685), .ZN(net_971), .A2(net_969) );
NAND2_X2 inst_1085 ( .A2(net_2023), .A1(net_1581), .ZN(net_432) );
INV_X2 inst_2328 ( .ZN(net_1012), .A(net_1011) );
NAND2_X2 inst_1667 ( .ZN(net_2692), .A2(net_1958), .A1(net_329) );
NAND2_X2 inst_1349 ( .A2(net_2328), .ZN(net_1091), .A1(net_617) );
DFFR_X1 inst_2655 ( .D(net_1502), .CK(net_2839), .RN(x2480), .Q(x434) );
NAND2_X1 inst_1720 ( .ZN(net_1612), .A1(net_752), .A2(net_695) );
OAI21_X2 inst_160 ( .ZN(net_2005), .B2(net_2004), .A(net_1714), .B1(net_419) );
NOR2_X2 inst_462 ( .ZN(net_2082), .A2(net_2081), .A1(net_975) );
NAND2_X4 inst_869 ( .A2(net_2603), .A1(net_2241), .ZN(net_1744) );
CLKBUF_X2 inst_3357 ( .A(net_3314), .Z(net_3315) );
DFFR_X1 inst_2646 ( .D(net_1479), .CK(net_3385), .RN(x2480), .Q(x339) );
OAI22_X4 inst_19 ( .A2(net_2782), .ZN(net_2102), .A1(net_634), .B1(net_133), .B2(net_39) );
OR2_X2 inst_8 ( .A2(net_2796), .A1(net_1826), .ZN(net_847) );
CLKBUF_X2 inst_2912 ( .A(net_2869), .Z(net_2870) );
NOR2_X2 inst_370 ( .A1(net_1997), .ZN(net_750), .A2(net_388) );
NAND2_X4 inst_762 ( .ZN(net_860), .A2(net_504), .A1(net_424) );
CLKBUF_X2 inst_3025 ( .A(net_2982), .Z(net_2983) );
INV_X2 inst_2224 ( .ZN(net_383), .A(net_360) );
NAND2_X2 inst_1265 ( .A1(net_1417), .A2(net_1232), .ZN(net_761) );
INV_X4 inst_2090 ( .ZN(net_1703), .A(net_1702) );
NAND2_X4 inst_965 ( .A1(net_2381), .ZN(net_2294), .A2(net_1954) );
CLKBUF_X2 inst_3267 ( .A(net_3224), .Z(net_3225) );
CLKBUF_X2 inst_3205 ( .A(net_3162), .Z(net_3163) );
NAND2_X1 inst_1686 ( .A1(net_778), .A2(net_686), .ZN(net_492) );
CLKBUF_X2 inst_3370 ( .A(net_2902), .Z(net_3328) );
INV_X4 inst_1914 ( .A(net_2383), .ZN(net_266) );
INV_X4 inst_1975 ( .A(net_1298), .ZN(net_786) );
INV_X4 inst_1890 ( .A(net_421), .ZN(net_364) );
INV_X2 inst_2308 ( .ZN(net_774), .A(net_204) );
NAND3_X2 inst_612 ( .A2(net_2585), .ZN(net_1160), .A3(net_1159), .A1(net_850) );
CLKBUF_X2 inst_2879 ( .A(net_2836), .Z(net_2837) );
INV_X8 inst_1789 ( .ZN(net_1787), .A(net_1786) );
NAND2_X1 inst_1692 ( .A2(net_2561), .A1(net_1934), .ZN(net_351) );
NAND2_X2 inst_1321 ( .A1(net_2711), .A2(net_2239), .ZN(net_965) );
NAND2_X4 inst_1012 ( .A2(net_2654), .A1(net_2652), .ZN(net_2557) );
NAND2_X4 inst_901 ( .ZN(net_1946), .A1(net_1102), .A2(net_330) );
INV_X2 inst_2338 ( .A(net_2358), .ZN(net_1263) );
INV_X4 inst_1956 ( .ZN(net_683), .A(net_682) );
CLKBUF_X2 inst_3017 ( .A(net_2974), .Z(net_2975) );
CLKBUF_X2 inst_3441 ( .A(net_3256), .Z(net_3399) );
NAND2_X4 inst_751 ( .A2(net_2239), .ZN(net_747), .A1(net_247) );
NAND2_X4 inst_845 ( .A2(net_2237), .ZN(net_1620), .A1(net_927) );
INV_X1 inst_2455 ( .A(net_2318), .ZN(net_601) );
CLKBUF_X2 inst_3149 ( .A(net_3106), .Z(net_3107) );
NAND2_X2 inst_1367 ( .A1(net_1189), .ZN(net_1172), .A2(net_813) );
INV_X1 inst_2471 ( .ZN(net_2281), .A(net_2280) );
INV_X2 inst_2403 ( .ZN(net_2594), .A(net_2593) );
NOR2_X2 inst_377 ( .A1(net_2551), .A2(net_1717), .ZN(net_806) );
INV_X4 inst_1934 ( .A(net_2102), .ZN(net_315) );
CLKBUF_X2 inst_3244 ( .A(net_3201), .Z(net_3202) );
CLKBUF_X2 inst_3098 ( .A(net_3055), .Z(net_3056) );
INV_X4 inst_2016 ( .A(net_1137), .ZN(net_1026) );
CLKBUF_X2 inst_3018 ( .A(net_2826), .Z(net_2976) );
CLKBUF_X2 inst_3078 ( .A(net_2948), .Z(net_3036) );
INV_X2 inst_2287 ( .ZN(net_40), .A(x831) );
NAND2_X2 inst_1460 ( .ZN(net_1621), .A2(net_1410), .A1(net_736) );
NAND2_X2 inst_1344 ( .A2(net_2249), .A1(net_1580), .ZN(net_1057) );
NAND2_X4 inst_885 ( .ZN(net_1851), .A1(net_1406), .A2(net_1022) );
DFFR_X1 inst_2630 ( .Q(net_2754), .D(net_2379), .CK(net_3087), .RN(x2480) );
CLKBUF_X2 inst_3053 ( .A(net_2982), .Z(net_3011) );
NAND2_X2 inst_1443 ( .ZN(net_1544), .A2(net_525), .A1(net_455) );
INV_X4 inst_2097 ( .ZN(net_1768), .A(net_1767) );
NAND2_X4 inst_928 ( .A2(net_2400), .ZN(net_2091), .A1(net_471) );
NAND2_X4 inst_1028 ( .ZN(net_2680), .A2(net_2679), .A1(net_2678) );
OAI21_X2 inst_107 ( .B1(net_1681), .ZN(net_552), .A(net_549), .B2(net_417) );
NOR2_X2 inst_393 ( .A2(net_1426), .A1(net_1223), .ZN(net_960) );
INV_X4 inst_2117 ( .ZN(net_1956), .A(net_1955) );
NAND2_X4 inst_990 ( .ZN(net_2435), .A1(net_2434), .A2(net_315) );
CLKBUF_X2 inst_3140 ( .A(net_3097), .Z(net_3098) );
CLKBUF_X2 inst_2999 ( .A(net_2898), .Z(net_2957) );
DFFR_X1 inst_2662 ( .D(net_1530), .CK(net_2893), .RN(x2480), .Q(x421) );
NAND2_X2 inst_1539 ( .A1(net_2483), .A2(net_2067), .ZN(net_2009) );
INV_X8 inst_1813 ( .A(net_2693), .ZN(net_2153) );
OAI21_X4 inst_92 ( .ZN(net_2199), .A(net_1831), .B2(net_237), .B1(net_155) );
NOR2_X2 inst_345 ( .A1(net_2297), .ZN(net_422), .A2(net_421) );
NAND2_X2 inst_1271 ( .A2(net_2323), .ZN(net_776), .A1(net_619) );
CLKBUF_X2 inst_3103 ( .A(net_3060), .Z(net_3061) );
NAND2_X1 inst_1718 ( .A1(net_2433), .A2(net_1964), .ZN(net_1203) );
NAND2_X2 inst_1050 ( .A2(net_1720), .ZN(net_547), .A1(net_516) );
INV_X2 inst_2366 ( .ZN(net_1742), .A(net_1219) );
INV_X2 inst_2321 ( .ZN(net_912), .A(net_911) );
CLKBUF_X2 inst_3304 ( .A(net_3261), .Z(net_3262) );
CLKBUF_X2 inst_3316 ( .A(net_3273), .Z(net_3274) );
NAND2_X2 inst_1296 ( .A2(net_2237), .ZN(net_893), .A1(net_892) );
INV_X4 inst_1852 ( .A(net_1245), .ZN(net_544) );
NOR3_X4 inst_200 ( .ZN(net_2670), .A3(net_2669), .A2(net_2666), .A1(net_2185) );
CLKBUF_X2 inst_3282 ( .A(net_3239), .Z(net_3240) );
OAI21_X4 inst_57 ( .B1(net_1585), .ZN(net_645), .A(net_644), .B2(net_37) );
NAND2_X2 inst_1557 ( .ZN(net_2117), .A2(net_2116), .A1(net_2115) );
INV_X8 inst_1750 ( .A(net_1826), .ZN(net_137) );
INV_X2 inst_2399 ( .ZN(net_2559), .A(net_347) );
INV_X2 inst_2236 ( .ZN(net_285), .A(net_158) );
CLKBUF_X2 inst_3368 ( .A(net_2855), .Z(net_3326) );
AOI22_X4 inst_2698 ( .ZN(net_2656), .A1(net_2655), .A2(net_2237), .B2(net_1689), .B1(net_1076) );
CLKBUF_X2 inst_3412 ( .A(net_3369), .Z(net_3370) );
NAND2_X2 inst_1553 ( .ZN(net_2100), .A2(net_1295), .A1(net_550) );
NAND2_X2 inst_1237 ( .ZN(net_2047), .A1(net_622), .A2(net_586) );
CLKBUF_X2 inst_3460 ( .A(net_3417), .Z(net_3418) );
DFFR_X2 inst_2518 ( .D(net_2281), .Q(net_1475), .CK(net_2817), .RN(x2480) );
AND2_X2 inst_2843 ( .ZN(net_1100), .A1(net_1099), .A2(net_918) );
INV_X4 inst_1888 ( .A(net_1104), .ZN(net_475) );
CLKBUF_X2 inst_3379 ( .A(net_3114), .Z(net_3337) );
INV_X8 inst_1763 ( .A(net_1087), .ZN(net_769) );
NAND2_X2 inst_1635 ( .ZN(net_2544), .A1(net_2352), .A2(net_2295) );
NAND2_X2 inst_1616 ( .ZN(net_2429), .A2(net_1677), .A1(net_1676) );
NAND2_X2 inst_1307 ( .ZN(net_921), .A2(net_523), .A1(net_458) );
CLKBUF_X2 inst_3310 ( .A(net_2970), .Z(net_3268) );
CLKBUF_X2 inst_3062 ( .A(net_3019), .Z(net_3020) );
INV_X4 inst_2075 ( .ZN(net_1591), .A(net_1590) );
INV_X4 inst_1911 ( .ZN(net_267), .A(net_257) );
NAND2_X2 inst_1500 ( .A1(net_1934), .A2(net_1851), .ZN(net_1813) );
AOI21_X2 inst_2805 ( .A(net_2602), .B1(net_2509), .B2(net_2409), .ZN(net_1278) );
INV_X8 inst_1825 ( .ZN(net_2383), .A(net_2382) );
NAND2_X2 inst_1094 ( .A2(net_2442), .A1(net_1352), .ZN(net_374) );
AND2_X2 inst_2851 ( .ZN(net_2741), .A1(net_2404), .A2(net_344) );
NAND2_X2 inst_1606 ( .ZN(net_2367), .A2(net_721), .A1(net_212) );
NAND3_X2 inst_585 ( .A3(net_1729), .A1(net_1609), .ZN(net_468), .A2(net_406) );
CLKBUF_X2 inst_2932 ( .A(net_2810), .Z(net_2890) );
NAND2_X4 inst_893 ( .A1(net_2008), .ZN(net_1888), .A2(net_908) );
NOR2_X2 inst_410 ( .ZN(net_1184), .A2(net_925), .A1(net_924) );
NOR2_X4 inst_316 ( .ZN(net_2476), .A1(net_2314), .A2(net_858) );
CLKBUF_X2 inst_3048 ( .A(net_3005), .Z(net_3006) );
NAND2_X1 inst_1699 ( .A2(net_1564), .ZN(net_192), .A1(net_187) );
NAND2_X4 inst_851 ( .ZN(net_1665), .A2(net_1664), .A1(net_1240) );
NAND2_X4 inst_831 ( .A2(net_2735), .A1(net_2734), .ZN(net_1509) );
NAND2_X2 inst_1174 ( .ZN(net_102), .A1(net_86), .A2(x701) );
NOR2_X2 inst_383 ( .A1(net_2466), .A2(net_1169), .ZN(net_899) );
NAND2_X4 inst_1023 ( .ZN(net_2635), .A1(net_2615), .A2(net_364) );
INV_X16 inst_2428 ( .A(net_2385), .ZN(net_2236) );
OAI21_X4 inst_50 ( .B1(net_1585), .A(net_651), .ZN(net_616), .B2(net_38) );
CLKBUF_X2 inst_3346 ( .A(net_3303), .Z(net_3304) );
NAND3_X4 inst_569 ( .ZN(net_1229), .A3(net_1228), .A1(net_1226), .A2(net_286) );
CLKBUF_X2 inst_2992 ( .A(net_2949), .Z(net_2950) );
CLKBUF_X2 inst_3186 ( .A(net_3143), .Z(net_3144) );
DFFR_X1 inst_2589 ( .Q(net_2759), .D(net_1185), .CK(net_3308), .RN(x2480) );
NAND2_X2 inst_1080 ( .A2(net_2536), .A1(net_488), .ZN(net_458) );
INV_X2 inst_2374 ( .ZN(net_1825), .A(net_98) );
NAND2_X2 inst_1124 ( .A1(net_619), .A2(net_242), .ZN(net_214) );
NAND3_X2 inst_678 ( .ZN(net_2449), .A3(net_2448), .A1(net_2446), .A2(net_1315) );
NAND2_X2 inst_1103 ( .A2(net_848), .ZN(net_565), .A1(net_312) );
CLKBUF_X2 inst_3259 ( .A(net_3114), .Z(net_3217) );
NAND2_X4 inst_854 ( .ZN(net_1671), .A2(net_764), .A1(net_572) );
CLKBUF_X2 inst_3375 ( .A(net_3332), .Z(net_3333) );
DFFR_X1 inst_2555 ( .QN(net_2787), .Q(net_1530), .D(net_886), .CK(net_3021), .RN(x2480) );
NAND2_X2 inst_1650 ( .ZN(net_2602), .A2(net_2601), .A1(net_2433) );
NAND4_X2 inst_549 ( .ZN(net_2364), .A3(net_2208), .A1(net_1727), .A4(net_1392), .A2(net_1257) );
NOR2_X4 inst_234 ( .ZN(net_1053), .A2(net_709), .A1(net_513) );
NAND2_X2 inst_1497 ( .ZN(net_1794), .A2(net_1653), .A1(net_1314) );
NAND4_X2 inst_522 ( .A3(net_1661), .A2(net_1340), .ZN(net_1253), .A1(net_1252), .A4(net_811) );
CLKBUF_X2 inst_2872 ( .A(net_2829), .Z(net_2830) );
NAND2_X4 inst_1002 ( .A1(net_2711), .ZN(net_2495), .A2(net_158) );
AOI21_X2 inst_2809 ( .B1(net_2428), .ZN(net_1451), .A(net_685), .B2(net_423) );
INV_X4 inst_1946 ( .ZN(net_117), .A(net_86) );
NOR2_X2 inst_478 ( .ZN(net_2536), .A2(net_2525), .A1(net_525) );
CLKBUF_X2 inst_3429 ( .A(net_3386), .Z(net_3387) );
CLKBUF_X2 inst_3380 ( .A(net_3251), .Z(net_3338) );
NAND2_X2 inst_1304 ( .A1(net_1778), .ZN(net_911), .A2(net_742) );
CLKBUF_X2 inst_3457 ( .A(net_3414), .Z(net_3415) );
NAND2_X2 inst_1328 ( .A1(net_2535), .ZN(net_984), .A2(net_981) );
NAND2_X2 inst_1618 ( .ZN(net_2451), .A2(net_2450), .A1(net_2449) );
NAND3_X2 inst_688 ( .ZN(net_2637), .A3(net_2636), .A1(net_2635), .A2(net_1337) );
CLKBUF_X2 inst_3292 ( .A(net_3044), .Z(net_3250) );
DFFR_X1 inst_2549 ( .QN(net_2794), .D(net_2720), .Q(net_1468), .CK(net_3425), .RN(x2480) );
INV_X4 inst_2126 ( .ZN(net_2010), .A(net_2009) );
INV_X8 inst_1749 ( .A(net_2132), .ZN(net_180) );
INV_X8 inst_1776 ( .ZN(net_1332), .A(net_1331) );
NAND2_X4 inst_804 ( .ZN(net_1260), .A2(net_1259), .A1(net_127) );
INV_X2 inst_2335 ( .ZN(net_1195), .A(net_276) );
CLKBUF_X2 inst_3290 ( .A(net_3247), .Z(net_3248) );
INV_X2 inst_2387 ( .ZN(net_2681), .A(net_2207) );
OR2_X2 inst_13 ( .A1(net_2740), .ZN(net_2436), .A2(net_987) );
NAND2_X4 inst_919 ( .ZN(net_2030), .A2(net_733), .A1(net_732) );
DFFR_X1 inst_2584 ( .D(net_2777), .CK(net_3330), .RN(x2480), .Q(x185) );
AOI21_X4 inst_2765 ( .A(net_2399), .B2(net_2396), .ZN(net_1056), .B1(net_1027) );
NAND3_X2 inst_598 ( .A3(net_2022), .ZN(net_851), .A2(net_731), .A1(net_432) );
CLKBUF_X2 inst_3156 ( .A(net_2949), .Z(net_3114) );
INV_X4 inst_1916 ( .ZN(net_283), .A(net_278) );
NAND2_X4 inst_799 ( .ZN(net_1237), .A2(net_1045), .A1(net_944) );
AOI22_X2 inst_2747 ( .A2(net_2754), .ZN(net_2552), .B1(net_296), .A1(net_284), .B2(x1808) );
NOR2_X4 inst_219 ( .A2(net_2562), .ZN(net_682), .A1(net_679) );
NAND2_X4 inst_738 ( .A1(net_1585), .A2(net_1496), .ZN(net_615) );
NAND2_X2 inst_1624 ( .ZN(net_2485), .A1(net_2481), .A2(net_1738) );
NAND2_X4 inst_719 ( .ZN(net_227), .A1(net_110), .A2(net_87) );
NAND2_X4 inst_840 ( .A1(net_2597), .ZN(net_1593), .A2(net_180) );
NAND2_X2 inst_1220 ( .A1(net_1585), .A2(net_1482), .ZN(net_636) );
AOI222_X1 inst_2755 ( .B1(net_2386), .C1(net_1943), .C2(net_1448), .A1(net_892), .A2(net_736), .ZN(net_289), .B2(net_209) );
INV_X4 inst_2181 ( .ZN(net_2565), .A(net_2564) );
NAND2_X2 inst_1456 ( .A2(net_1702), .ZN(net_1609), .A1(net_405) );
INV_X8 inst_1819 ( .ZN(net_2287), .A(net_2286) );
INV_X8 inst_1797 ( .A(net_1908), .ZN(net_1905) );
NOR2_X4 inst_255 ( .A2(net_1672), .ZN(net_1393), .A1(net_494) );
AOI22_X2 inst_2726 ( .A2(net_2769), .ZN(net_1274), .B1(net_296), .A1(net_283), .B2(x1620) );
NOR2_X2 inst_453 ( .ZN(net_1997), .A1(net_1994), .A2(net_1509) );
CLKBUF_X2 inst_3167 ( .A(net_3124), .Z(net_3125) );
NAND2_X2 inst_1134 ( .A2(net_243), .ZN(net_197), .A1(net_158) );
NOR2_X1 inst_493 ( .A2(net_2788), .ZN(net_925), .A1(net_634) );
INV_X2 inst_2204 ( .A(net_2461), .ZN(net_497) );
OAI22_X2 inst_23 ( .B2(net_2797), .B1(net_633), .ZN(net_182), .A1(net_143), .A2(net_60) );
AOI22_X2 inst_2708 ( .A2(net_2778), .ZN(net_299), .A1(net_295), .B1(net_126), .B2(x1719) );
NAND2_X2 inst_1113 ( .A2(net_586), .ZN(net_566), .A1(net_247) );
INV_X8 inst_1822 ( .ZN(net_2320), .A(net_2319) );
NAND2_X2 inst_1609 ( .ZN(net_2387), .A2(net_2386), .A1(net_2384) );
NOR2_X2 inst_408 ( .A1(net_2401), .ZN(net_1169), .A2(net_343) );
DFFR_X1 inst_2592 ( .D(net_2765), .CK(net_3150), .RN(x2480), .Q(x451) );
NAND2_X2 inst_1144 ( .A2(net_2328), .A1(net_203), .ZN(net_183) );
NOR2_X4 inst_325 ( .ZN(net_2609), .A2(net_2608), .A1(net_2607) );
NAND2_X4 inst_812 ( .A1(net_2727), .A2(net_1439), .ZN(net_1323) );
CLKBUF_X2 inst_3116 ( .A(net_3073), .Z(net_3074) );
DFFR_X1 inst_2568 ( .D(net_2776), .CK(net_3249), .RN(x2480), .Q(x128) );
NAND2_X2 inst_1197 ( .A1(net_1585), .A2(net_1516), .ZN(net_588) );
INV_X2 inst_2295 ( .ZN(net_33), .A(x562) );
OAI21_X2 inst_179 ( .ZN(net_2661), .B2(net_2660), .B1(net_1887), .A(net_316) );
NAND2_X4 inst_955 ( .ZN(net_2240), .A2(net_1283), .A1(net_1282) );
NAND2_X1 inst_1730 ( .ZN(net_2612), .A1(net_2610), .A2(net_2435) );
OAI21_X2 inst_114 ( .A(net_1380), .B2(net_319), .ZN(net_259), .B1(net_255) );
INV_X2 inst_2278 ( .ZN(net_49), .A(x2049) );
CLKBUF_X2 inst_3028 ( .A(net_2985), .Z(net_2986) );
INV_X4 inst_2191 ( .ZN(net_2668), .A(net_2667) );
OAI21_X4 inst_76 ( .ZN(net_1731), .B1(net_1585), .A(net_636), .B2(net_56) );
NAND3_X2 inst_617 ( .A3(net_1440), .ZN(net_1289), .A1(net_379), .A2(net_353) );
NAND2_X2 inst_1127 ( .A1(net_234), .A2(net_227), .ZN(net_208) );
OAI21_X2 inst_172 ( .ZN(net_2391), .B2(net_2390), .B1(net_2389), .A(net_2388) );
NOR2_X2 inst_362 ( .A1(net_1008), .ZN(net_218), .A2(net_142) );
NAND2_X2 inst_1530 ( .A1(net_2657), .ZN(net_1981), .A2(net_1980) );
NOR2_X4 inst_277 ( .A1(net_2396), .A2(net_1917), .ZN(net_1814) );
NAND2_X2 inst_1510 ( .ZN(net_1871), .A1(net_1870), .A2(net_1085) );
OAI21_X4 inst_83 ( .ZN(net_1937), .B2(net_156), .A(net_111), .B1(net_61) );
OAI21_X2 inst_121 ( .B2(net_2551), .B1(net_1416), .ZN(net_702), .A(net_549) );
NOR2_X4 inst_306 ( .ZN(net_2300), .A2(net_2090), .A1(net_2089) );
NAND4_X2 inst_534 ( .A4(net_1846), .ZN(net_1774), .A3(net_1773), .A2(net_1772), .A1(net_1771) );
NAND2_X2 inst_1065 ( .A1(net_729), .ZN(net_494), .A2(net_493) );
NAND2_X2 inst_1057 ( .A2(net_1362), .ZN(net_523), .A1(net_522) );
CLKBUF_X2 inst_3386 ( .A(net_3343), .Z(net_3344) );
CLKBUF_X2 inst_3095 ( .A(net_3052), .Z(net_3053) );
NAND2_X1 inst_1715 ( .A1(net_1906), .ZN(net_986), .A2(net_980) );
OAI21_X2 inst_140 ( .B2(net_1910), .B1(net_1906), .ZN(net_1306), .A(net_1305) );
NOR2_X4 inst_267 ( .A1(net_2174), .ZN(net_1599), .A2(net_1574) );
AND2_X2 inst_2842 ( .A1(net_1914), .ZN(net_1078), .A2(net_1077) );
AND3_X4 inst_2824 ( .ZN(net_2180), .A1(net_1597), .A2(net_1249), .A3(net_95) );
AND2_X4 inst_2836 ( .ZN(net_2212), .A2(net_2211), .A1(net_2210) );
INV_X4 inst_2084 ( .A(net_1859), .ZN(net_1653) );
NAND2_X4 inst_748 ( .A2(net_2111), .A1(net_1194), .ZN(net_728) );
AND2_X4 inst_2839 ( .ZN(net_2653), .A2(net_1136), .A1(net_893) );
NAND2_X4 inst_716 ( .A2(net_1943), .ZN(net_666), .A1(net_173) );
AOI21_X4 inst_2770 ( .A(net_1915), .B2(net_1817), .ZN(net_1550), .B1(net_1549) );
INV_X4 inst_1906 ( .A(net_2046), .ZN(net_311) );
NAND4_X2 inst_530 ( .A3(net_2263), .A2(net_1778), .ZN(net_1642), .A4(net_742), .A1(net_610) );
NAND2_X4 inst_792 ( .A2(net_2505), .ZN(net_1179), .A1(net_387) );
INV_X4 inst_2024 ( .A(net_1604), .ZN(net_1102) );
CLKBUF_X2 inst_3124 ( .A(net_2962), .Z(net_3082) );
CLKBUF_X2 inst_3444 ( .A(net_3401), .Z(net_3402) );
CLKBUF_X2 inst_2952 ( .A(net_2909), .Z(net_2910) );
NAND2_X2 inst_1353 ( .A1(net_2579), .ZN(net_1105), .A2(net_991) );
DFFR_X2 inst_2502 ( .D(net_1878), .Q(net_1473), .CK(net_2885), .RN(x2480) );
NAND2_X4 inst_803 ( .A2(net_2420), .ZN(net_1249), .A1(net_941) );
CLKBUF_X2 inst_2909 ( .A(net_2835), .Z(net_2867) );
INV_X4 inst_1986 ( .A(net_2070), .ZN(net_833) );
INV_X4 inst_1949 ( .ZN(net_2014), .A(net_681) );
INV_X2 inst_2216 ( .A(net_2071), .ZN(net_449) );
NAND2_X4 inst_769 ( .ZN(net_1908), .A1(net_699), .A2(net_331) );
OAI21_X2 inst_174 ( .B2(net_2596), .ZN(net_2556), .B1(net_2553), .A(net_2552) );
CLKBUF_X2 inst_3135 ( .A(net_3092), .Z(net_3093) );
INV_X2 inst_2348 ( .ZN(net_2438), .A(net_1998) );
NAND2_X2 inst_1200 ( .A1(net_1585), .A2(net_1503), .ZN(net_592) );
CLKBUF_X2 inst_2988 ( .A(net_2945), .Z(net_2946) );
NAND3_X2 inst_662 ( .ZN(net_2127), .A3(net_2126), .A2(net_2125), .A1(net_2124) );
NAND3_X1 inst_701 ( .A1(net_2165), .ZN(net_1161), .A3(net_1159), .A2(net_867) );
CLKBUF_X2 inst_2911 ( .A(net_2868), .Z(net_2869) );
INV_X2 inst_2380 ( .A(net_1918), .ZN(net_1917) );
NAND2_X2 inst_1533 ( .ZN(net_1991), .A2(net_1990), .A1(net_454) );
INV_X4 inst_2105 ( .ZN(net_1832), .A(net_1224) );
NAND2_X2 inst_1199 ( .A1(net_1585), .A2(net_1483), .ZN(net_590) );
OR2_X4 inst_5 ( .A2(net_1652), .ZN(net_1511), .A1(net_426) );
CLKBUF_X2 inst_3021 ( .A(net_2978), .Z(net_2979) );
NAND2_X4 inst_729 ( .A2(net_1515), .ZN(net_122), .A1(net_121) );
INV_X4 inst_2157 ( .A(net_2680), .ZN(net_2356) );
NAND2_X2 inst_1662 ( .ZN(net_2658), .A2(net_1859), .A1(net_1856) );
AOI21_X2 inst_2783 ( .ZN(net_2684), .B2(net_1265), .B1(net_1154), .A(net_999) );
INV_X4 inst_1859 ( .A(net_1718), .ZN(net_433) );
NOR2_X4 inst_213 ( .A1(net_2453), .A2(net_1905), .ZN(net_488) );
NAND2_X2 inst_1465 ( .ZN(net_1634), .A1(net_1633), .A2(net_282) );
NAND3_X2 inst_604 ( .A2(net_2351), .A3(net_1927), .ZN(net_951), .A1(net_948) );
OAI21_X4 inst_53 ( .B1(net_1585), .ZN(net_621), .A(net_620), .B2(net_58) );
AOI21_X2 inst_2815 ( .ZN(net_2257), .B1(net_2256), .A(net_766), .B2(net_613) );
NAND2_X4 inst_1007 ( .ZN(net_2530), .A2(net_2525), .A1(net_1545) );
NOR3_X2 inst_205 ( .A3(net_2329), .A1(net_1843), .ZN(net_1372), .A2(net_1371) );
NAND2_X2 inst_1645 ( .ZN(net_2590), .A1(net_2589), .A2(net_187) );
NAND2_X2 inst_1285 ( .A2(net_2506), .A1(net_1991), .ZN(net_1215) );
NOR2_X2 inst_380 ( .A1(net_1579), .A2(net_934), .ZN(net_818) );
NAND2_X2 inst_1179 ( .ZN(net_91), .A1(net_86), .A2(x651) );
CLKBUF_X2 inst_3337 ( .A(net_3294), .Z(net_3295) );
DFFR_X1 inst_2614 ( .Q(net_2769), .D(net_813), .CK(net_3010), .RN(x2480) );
NAND3_X2 inst_651 ( .A3(net_2379), .ZN(net_1954), .A1(net_1891), .A2(net_939) );
NOR2_X4 inst_292 ( .ZN(net_2128), .A2(net_1698), .A1(net_1697) );
NAND2_X4 inst_999 ( .ZN(net_2477), .A1(net_2476), .A2(net_552) );
CLKBUF_X2 inst_2883 ( .A(net_2827), .Z(net_2841) );
INV_X4 inst_2111 ( .A(net_1911), .ZN(net_1910) );
INV_X4 inst_2012 ( .A(net_1051), .ZN(net_1010) );
INV_X8 inst_1846 ( .ZN(net_2592), .A(net_2589) );
NAND2_X2 inst_1157 ( .ZN(net_124), .A1(net_112), .A2(net_74) );
INV_X4 inst_2139 ( .ZN(net_2171), .A(net_2170) );
NAND2_X2 inst_1515 ( .ZN(net_1885), .A1(net_1884), .A2(net_317) );
NAND2_X2 inst_1463 ( .ZN(net_1629), .A1(net_1628), .A2(net_1094) );
OAI211_X2 inst_186 ( .C1(net_2549), .C2(net_1231), .A(net_1175), .B(net_952), .ZN(net_858) );
NAND2_X4 inst_706 ( .A2(net_570), .ZN(net_510), .A1(net_463) );
NAND2_X4 inst_759 ( .ZN(net_825), .A2(net_654), .A1(net_653) );
CLKBUF_X2 inst_3071 ( .A(net_3028), .Z(net_3029) );
INV_X8 inst_1782 ( .ZN(net_1547), .A(net_1546) );
INV_X4 inst_2061 ( .ZN(net_1384), .A(net_1383) );
CLKBUF_X2 inst_2951 ( .A(net_2861), .Z(net_2909) );
NAND2_X4 inst_863 ( .ZN(net_1704), .A1(net_713), .A2(net_250) );
NAND2_X4 inst_839 ( .A2(net_2530), .ZN(net_1583), .A1(net_772) );
NAND2_X4 inst_1015 ( .ZN(net_2588), .A2(net_2587), .A1(net_2585) );
NAND2_X2 inst_1472 ( .A2(net_2133), .ZN(net_1692), .A1(net_1688) );
NOR2_X4 inst_240 ( .A1(net_2689), .A2(net_1182), .ZN(net_1139) );
NAND2_X2 inst_1385 ( .ZN(net_1259), .A1(net_1258), .A2(x761) );
OAI21_X2 inst_110 ( .A(net_1388), .B2(net_571), .ZN(net_513), .B1(net_508) );
NAND2_X2 inst_1573 ( .ZN(net_2170), .A1(net_705), .A2(net_704) );
NAND2_X2 inst_1183 ( .ZN(net_88), .A1(net_86), .A2(x899) );
NAND2_X2 inst_1390 ( .ZN(net_1277), .A2(net_1275), .A1(net_1036) );
INV_X4 inst_2047 ( .A(net_2198), .ZN(net_1252) );
CLKBUF_X2 inst_3213 ( .A(net_3170), .Z(net_3171) );
NOR2_X4 inst_229 ( .A2(net_2288), .ZN(net_969), .A1(net_367) );
DFFR_X1 inst_2535 ( .QN(net_2797), .D(net_1754), .Q(net_1476), .CK(net_3280), .RN(x2480) );
OAI21_X4 inst_99 ( .ZN(net_2450), .B1(net_2445), .B2(net_1967), .A(net_1966) );
INV_X2 inst_2282 ( .ZN(net_45), .A(x1868) );
NAND2_X2 inst_1489 ( .ZN(net_1743), .A1(net_1220), .A2(net_1218) );
INV_X16 inst_2415 ( .A(net_1240), .ZN(net_1069) );
NAND2_X2 inst_1661 ( .ZN(net_2649), .A1(net_1839), .A2(net_893) );
CLKBUF_X2 inst_3288 ( .A(net_3245), .Z(net_3246) );
INV_X2 inst_2262 ( .ZN(net_65), .A(x1710) );
INV_X4 inst_2059 ( .ZN(net_1362), .A(net_1359) );
CLKBUF_X2 inst_2949 ( .A(net_2827), .Z(net_2907) );
INV_X16 inst_2414 ( .A(net_2182), .ZN(net_1007) );
NAND2_X2 inst_1394 ( .A2(net_1547), .ZN(net_1294), .A1(net_461) );
NAND2_X2 inst_1160 ( .A1(net_133), .ZN(net_120), .A2(net_77) );
INV_X4 inst_2131 ( .ZN(net_2096), .A(net_2095) );
NOR2_X4 inst_283 ( .ZN(net_1953), .A2(net_857), .A1(net_237) );
NOR2_X4 inst_311 ( .ZN(net_2376), .A2(net_2072), .A1(net_2013) );
CLKBUF_X2 inst_3406 ( .A(net_3282), .Z(net_3364) );
DFFR_X2 inst_2519 ( .D(net_2058), .Q(net_1465), .CK(net_3183), .RN(x2480) );
INV_X8 inst_1808 ( .A(net_2179), .ZN(net_2112) );
NAND2_X2 inst_1597 ( .ZN(net_2312), .A2(net_1453), .A1(net_946) );
INV_X4 inst_1876 ( .A(net_2000), .ZN(net_456) );
NAND2_X4 inst_988 ( .ZN(net_2407), .A2(net_2229), .A1(net_1888) );
INV_X2 inst_2203 ( .A(net_2520), .ZN(net_507) );
OAI21_X2 inst_169 ( .ZN(net_2314), .B2(net_2313), .B1(net_2311), .A(net_2310) );
NOR2_X2 inst_421 ( .A1(net_2484), .A2(net_2071), .ZN(net_1354) );
NAND2_X2 inst_1315 ( .A2(net_2581), .ZN(net_953), .A1(net_469) );
NAND4_X2 inst_555 ( .ZN(net_2627), .A3(net_2625), .A4(net_1867), .A1(net_1396), .A2(net_1348) );
INV_X2 inst_2392 ( .ZN(net_2357), .A(net_2356) );
NAND2_X4 inst_816 ( .ZN(net_1912), .A2(net_1686), .A1(net_1445) );
NOR2_X2 inst_431 ( .ZN(net_1436), .A1(net_1360), .A2(net_438) );
AOI21_X2 inst_2798 ( .B1(net_2339), .A(net_1167), .ZN(net_1034), .B2(net_1032) );
NOR2_X2 inst_348 ( .A1(net_994), .ZN(net_396), .A2(net_357) );
INV_X4 inst_1930 ( .A(net_1008), .ZN(net_242) );
NAND2_X2 inst_1184 ( .ZN(net_653), .A1(net_86), .A2(x609) );
NAND2_X4 inst_889 ( .A2(net_2362), .ZN(net_1862), .A1(net_1720) );
NAND3_X4 inst_577 ( .ZN(net_2241), .A3(net_2240), .A1(net_1785), .A2(net_506) );
INV_X2 inst_2293 ( .ZN(net_35), .A(x574) );
INV_X2 inst_2379 ( .A(net_1912), .ZN(net_1909) );
NAND2_X2 inst_1364 ( .A2(net_1287), .A1(net_1180), .ZN(net_1156) );
NAND3_X2 inst_656 ( .ZN(net_2018), .A1(net_2017), .A2(net_1643), .A3(net_1312) );
CLKBUF_X2 inst_2865 ( .A(net_2810), .Z(net_2823) );
NAND3_X2 inst_645 ( .ZN(net_1864), .A3(net_1862), .A1(net_1724), .A2(net_1678) );
OAI21_X4 inst_45 ( .B2(net_2132), .ZN(net_256), .B1(net_255), .A(net_190) );
CLKBUF_X2 inst_3041 ( .A(net_2930), .Z(net_2999) );
NAND2_X2 inst_1108 ( .ZN(net_262), .A1(net_214), .A2(net_207) );
AOI22_X2 inst_2719 ( .A2(net_2777), .ZN(net_868), .A1(net_283), .B1(net_126), .B2(x1593) );
INV_X2 inst_2352 ( .A(net_2671), .ZN(net_1568) );
NOR2_X4 inst_269 ( .A2(net_2091), .ZN(net_1661), .A1(net_1402) );
CLKBUF_X2 inst_3093 ( .A(net_2861), .Z(net_3051) );
NAND2_X2 inst_1190 ( .A1(net_2386), .ZN(net_575), .A2(net_217) );
NOR2_X2 inst_458 ( .ZN(net_2069), .A1(net_2068), .A2(net_1610) );
NOR2_X2 inst_444 ( .ZN(net_1782), .A2(net_1288), .A1(net_454) );
NAND2_X2 inst_1562 ( .ZN(net_2125), .A1(net_1602), .A2(net_736) );
INV_X4 inst_1922 ( .A(net_330), .ZN(net_313) );
CLKBUF_X2 inst_3361 ( .A(net_3318), .Z(net_3319) );
CLKBUF_X2 inst_3170 ( .A(net_3127), .Z(net_3128) );
DFFR_X1 inst_2544 ( .D(net_1736), .Q(net_69), .CK(net_3083), .RN(x2480) );
NAND2_X4 inst_741 ( .A2(net_1632), .A1(net_1429), .ZN(net_672) );
CLKBUF_X2 inst_3232 ( .A(net_3189), .Z(net_3190) );
NAND4_X2 inst_514 ( .A1(net_2693), .A2(net_2585), .A4(net_2165), .A3(net_1158), .ZN(net_955) );
NAND2_X2 inst_1541 ( .ZN(net_2028), .A2(net_2025), .A1(net_2024) );
CLKBUF_X2 inst_3343 ( .A(net_3300), .Z(net_3301) );
NAND3_X2 inst_685 ( .ZN(net_2596), .A2(net_2593), .A3(net_2555), .A1(net_2554) );
NAND2_X2 inst_1350 ( .A2(net_2320), .A1(net_1191), .ZN(net_1092) );
OAI21_X4 inst_63 ( .ZN(net_977), .A(net_914), .B2(net_545), .B1(net_460) );
CLKBUF_X2 inst_3012 ( .A(net_2969), .Z(net_2970) );
DFFR_X1 inst_2635 ( .D(net_72), .CK(net_3337), .RN(x2480), .Q(x193) );
OAI21_X2 inst_119 ( .B1(net_1585), .ZN(net_643), .A(net_642), .B2(net_44) );
CLKBUF_X2 inst_3181 ( .A(net_3138), .Z(net_3139) );
NAND2_X4 inst_939 ( .ZN(net_2157), .A2(net_2060), .A1(net_1399) );
AND2_X4 inst_2828 ( .A1(net_2362), .A2(net_1720), .ZN(net_1510) );
NAND2_X2 inst_1543 ( .A2(net_2655), .ZN(net_2044), .A1(net_721) );
AOI21_X2 inst_2801 ( .A(net_2569), .B2(net_2390), .B1(net_1201), .ZN(net_1143) );
NAND2_X2 inst_1118 ( .A2(net_245), .A1(net_242), .ZN(net_224) );
INV_X2 inst_2303 ( .A(net_713), .ZN(net_712) );
CLKBUF_X2 inst_3363 ( .A(net_3320), .Z(net_3321) );
NAND2_X2 inst_1233 ( .A1(net_1585), .A2(net_1506), .ZN(net_651) );
CLKBUF_X2 inst_2924 ( .A(net_2881), .Z(net_2882) );
CLKBUF_X2 inst_3432 ( .A(net_3389), .Z(net_3390) );
NAND2_X4 inst_1019 ( .ZN(net_2601), .A1(net_1765), .A2(net_751) );
INV_X4 inst_2006 ( .ZN(net_973), .A(net_568) );
NOR2_X2 inst_473 ( .ZN(net_2389), .A1(net_1618), .A2(net_690) );
INV_X8 inst_1827 ( .ZN(net_2395), .A(net_2394) );
NAND2_X2 inst_1131 ( .A2(net_2237), .A1(net_244), .ZN(net_202) );
NAND2_X2 inst_1357 ( .ZN(net_1132), .A2(net_1131), .A1(net_738) );
NAND2_X4 inst_742 ( .A2(net_1725), .ZN(net_681), .A1(net_680) );
INV_X2 inst_2211 ( .A(net_1707), .ZN(net_413) );
NAND3_X2 inst_691 ( .ZN(net_2664), .A2(net_2663), .A1(net_1886), .A3(net_855) );
NOR2_X2 inst_427 ( .A2(net_2691), .A1(net_1876), .ZN(net_1403) );
DFFR_X1 inst_2619 ( .D(net_151), .CK(net_3163), .RN(x2480), .Q(x0) );
CLKBUF_X2 inst_3083 ( .A(net_3040), .Z(net_3041) );
NAND2_X1 inst_1695 ( .A2(net_1689), .A1(net_622), .ZN(net_251) );
CLKBUF_X2 inst_3465 ( .A(net_3422), .Z(net_3423) );
INV_X4 inst_2033 ( .A(net_2515), .ZN(net_1163) );
INV_X4 inst_2144 ( .ZN(net_2232), .A(net_990) );
NAND2_X4 inst_770 ( .A1(net_1332), .ZN(net_993), .A2(net_421) );
NAND3_X4 inst_565 ( .A2(net_740), .A1(net_600), .ZN(net_275), .A3(net_175) );
DFFR_X1 inst_2559 ( .QN(net_2788), .Q(net_1463), .D(net_1346), .CK(net_3054), .RN(x2480) );
INV_X4 inst_1971 ( .A(net_2258), .ZN(net_765) );
OAI21_X2 inst_138 ( .B2(net_1718), .B1(net_1454), .ZN(net_1153), .A(net_503) );
NAND3_X2 inst_622 ( .A3(net_2606), .ZN(net_1346), .A2(net_1345), .A1(net_1342) );
INV_X4 inst_1955 ( .A(net_670), .ZN(net_669) );
NAND2_X2 inst_1404 ( .A2(net_1714), .A1(net_1329), .ZN(net_1321) );
CLKBUF_X2 inst_2989 ( .A(net_2946), .Z(net_2947) );
AOI21_X2 inst_2810 ( .ZN(net_1809), .B2(net_995), .A(net_937), .B1(net_860) );
NOR2_X2 inst_409 ( .ZN(net_1178), .A2(net_1177), .A1(net_416) );
INV_X2 inst_2288 ( .ZN(net_39), .A(x1280) );
NAND2_X2 inst_1269 ( .ZN(net_777), .A2(net_776), .A1(net_775) );
NAND2_X2 inst_1339 ( .A1(net_1204), .ZN(net_1031), .A2(net_864) );
NAND2_X4 inst_899 ( .ZN(net_1942), .A2(net_1941), .A1(net_649) );
INV_X8 inst_1834 ( .ZN(net_2433), .A(net_2432) );
NOR2_X4 inst_312 ( .ZN(net_2385), .A2(net_1895), .A1(net_1894) );
NAND2_X4 inst_977 ( .ZN(net_2373), .A2(net_2372), .A1(net_2371) );
CLKBUF_X2 inst_3241 ( .A(net_2987), .Z(net_3199) );
AOI22_X2 inst_2704 ( .A2(net_2763), .ZN(net_297), .B1(net_296), .A1(net_284), .B2(x1863) );
INV_X2 inst_2228 ( .A(net_2398), .ZN(net_347) );
NAND2_X2 inst_1620 ( .ZN(net_2467), .A1(net_2464), .A2(net_1632) );
NOR2_X4 inst_309 ( .ZN(net_2315), .A2(net_1606), .A1(net_1605) );
CLKBUF_X2 inst_3416 ( .A(net_3373), .Z(net_3374) );
NOR2_X2 inst_347 ( .A2(net_2603), .A1(net_1288), .ZN(net_398) );
NAND2_X4 inst_768 ( .A2(net_1905), .ZN(net_981), .A1(net_980) );
NAND3_X2 inst_663 ( .A1(net_2671), .ZN(net_2184), .A3(net_2183), .A2(net_1164) );
INV_X4 inst_2121 ( .ZN(net_1985), .A(net_137) );
INV_X4 inst_2149 ( .A(net_2680), .ZN(net_2288) );
NOR2_X4 inst_297 ( .A2(net_2238), .ZN(net_2193), .A1(net_1317) );
NAND2_X4 inst_755 ( .ZN(net_785), .A2(net_203), .A1(net_158) );
CLKBUF_X2 inst_3227 ( .A(net_3184), .Z(net_3185) );
DFFR_X2 inst_2477 ( .Q(net_1529), .D(net_1378), .CK(net_2835), .RN(x2480) );
NAND2_X1 inst_1724 ( .A2(net_2321), .ZN(net_1709), .A1(net_180) );
NAND2_X2 inst_1395 ( .A2(net_1899), .A1(net_1547), .ZN(net_1295) );
CLKBUF_X2 inst_3436 ( .A(net_3322), .Z(net_3394) );
DFFR_X1 inst_2610 ( .D(net_2771), .CK(net_3413), .RN(x2480), .Q(x316) );
INV_X4 inst_2188 ( .ZN(net_2650), .A(net_2649) );
AOI22_X4 inst_2694 ( .A2(net_2538), .B1(net_2456), .A1(net_2184), .ZN(net_1791), .B2(net_529) );
CLKBUF_X2 inst_3351 ( .A(net_2954), .Z(net_3309) );
INV_X4 inst_1875 ( .A(net_527), .ZN(net_401) );
NAND2_X2 inst_1043 ( .A1(net_1444), .A2(net_1141), .ZN(net_562) );
INV_X4 inst_1867 ( .A(net_671), .ZN(net_484) );
CLKBUF_X2 inst_3190 ( .A(net_3147), .Z(net_3148) );
OAI21_X2 inst_162 ( .ZN(net_2066), .A(net_2064), .B2(net_2061), .B1(net_583) );
INV_X4 inst_1968 ( .A(net_2201), .ZN(net_754) );
CLKBUF_X2 inst_3308 ( .A(net_3265), .Z(net_3266) );
INV_X2 inst_2290 ( .ZN(net_38), .A(x638) );
INV_X8 inst_1792 ( .A(net_1982), .ZN(net_1824) );
CLKBUF_X2 inst_3397 ( .A(net_3354), .Z(net_3355) );
NAND2_X2 inst_1330 ( .ZN(net_988), .A1(net_616), .A2(net_180) );
CLKBUF_X2 inst_3353 ( .A(net_3310), .Z(net_3311) );
INV_X4 inst_1898 ( .A(net_2268), .ZN(net_359) );
AND2_X4 inst_2829 ( .ZN(net_1656), .A1(net_1235), .A2(net_1097) );
NAND2_X1 inst_1714 ( .A1(net_2277), .A2(net_1211), .ZN(net_906) );
CLKBUF_X2 inst_3342 ( .A(net_3299), .Z(net_3300) );
NAND2_X2 inst_1098 ( .A1(net_2562), .A2(net_809), .ZN(net_354) );
DFFR_X1 inst_2621 ( .Q(net_2762), .D(net_1120), .CK(net_3074), .RN(x2480) );
NAND2_X2 inst_1496 ( .A2(net_2711), .ZN(net_1781), .A1(net_586) );
INV_X16 inst_2443 ( .ZN(net_2587), .A(net_2586) );
NAND2_X2 inst_1565 ( .ZN(net_2146), .A1(net_2145), .A2(net_1020) );
NAND2_X4 inst_924 ( .A2(net_2062), .ZN(net_2054), .A1(net_1082) );
NOR2_X4 inst_303 ( .ZN(net_2256), .A2(net_966), .A1(net_963) );
NAND2_X4 inst_723 ( .A1(net_628), .ZN(net_247), .A2(net_103) );
NOR2_X4 inst_287 ( .ZN(net_2056), .A1(net_1132), .A2(net_238) );
INV_X16 inst_2444 ( .ZN(net_2603), .A(net_2601) );
NOR2_X2 inst_426 ( .A1(net_2255), .ZN(net_1391), .A2(net_1390) );
NAND3_X2 inst_618 ( .A3(net_2672), .A2(net_1923), .ZN(net_1308), .A1(net_1307) );
CLKBUF_X2 inst_3145 ( .A(net_2814), .Z(net_3103) );
DFFR_X1 inst_2577 ( .D(net_2751), .CK(net_3226), .RN(x2480), .Q(x114) );
CLKBUF_X2 inst_3263 ( .A(net_3009), .Z(net_3221) );
NAND2_X2 inst_1647 ( .ZN(net_2598), .A2(net_2597), .A1(net_2237) );
NAND3_X2 inst_648 ( .ZN(net_1930), .A1(net_1929), .A3(net_1845), .A2(net_1384) );
CLKBUF_X2 inst_3094 ( .A(net_3051), .Z(net_3052) );
CLKBUF_X2 inst_3057 ( .A(net_3014), .Z(net_3015) );
INV_X1 inst_2462 ( .ZN(net_1270), .A(net_1269) );
NAND2_X2 inst_1275 ( .ZN(net_793), .A2(net_736), .A1(net_245) );
CLKBUF_X2 inst_2903 ( .A(net_2860), .Z(net_2861) );
NOR2_X4 inst_270 ( .A2(net_2032), .ZN(net_1673), .A1(net_258) );
INV_X4 inst_1901 ( .A(net_1559), .ZN(net_384) );
NOR2_X2 inst_474 ( .A2(net_2804), .ZN(net_2420), .A1(net_2419) );
OAI22_X2 inst_26 ( .A2(net_2794), .ZN(net_928), .A1(net_634), .B1(net_112), .B2(net_66) );
INV_X4 inst_2067 ( .ZN(net_1514), .A(net_1513) );
NAND2_X4 inst_984 ( .A2(net_2562), .ZN(net_2392), .A1(net_352) );
NAND3_X2 inst_626 ( .A3(net_2728), .A1(net_2696), .A2(net_2286), .ZN(net_1899) );
CLKBUF_X2 inst_2882 ( .A(net_2833), .Z(net_2840) );
INV_X4 inst_2064 ( .ZN(net_1454), .A(net_1453) );
NAND2_X2 inst_1376 ( .A1(net_2275), .ZN(net_1211), .A2(net_866) );
AOI21_X4 inst_2777 ( .A(net_2396), .ZN(net_2207), .B1(net_1138), .B2(net_397) );
INV_X2 inst_2266 ( .ZN(net_61), .A(x1582) );
NAND2_X2 inst_1292 ( .ZN(net_881), .A1(net_880), .A2(net_307) );
DFFR_X1 inst_2552 ( .D(net_2703), .Q(net_76), .CK(net_3276), .RN(x2480) );
INV_X16 inst_2446 ( .ZN(net_2726), .A(net_2725) );
INV_X4 inst_1963 ( .A(net_997), .ZN(net_713) );
NAND3_X2 inst_631 ( .A1(net_2567), .A3(net_2129), .A2(net_2096), .ZN(net_1573) );
NAND2_X2 inst_1056 ( .A2(net_972), .A1(net_962), .ZN(net_526) );
NAND2_X2 inst_1659 ( .ZN(net_2643), .A1(net_2642), .A2(net_744) );
NAND2_X4 inst_798 ( .A1(net_1767), .ZN(net_1236), .A2(net_385) );
DFFR_X2 inst_2514 ( .D(net_1983), .Q(net_1474), .CK(net_2862), .RN(x2480) );
NOR2_X2 inst_398 ( .A2(net_1288), .ZN(net_1033), .A1(net_1032) );
NAND2_X2 inst_1128 ( .A1(net_1009), .ZN(net_206), .A2(net_200) );
NOR2_X2 inst_436 ( .A1(net_2274), .ZN(net_1608), .A2(net_1607) );
CLKBUF_X2 inst_3222 ( .A(net_2903), .Z(net_3180) );
NAND2_X2 inst_1434 ( .ZN(net_1412), .A1(net_1411), .A2(net_802) );
INV_X4 inst_1886 ( .ZN(net_525), .A(net_444) );
INV_X8 inst_1745 ( .A(net_2327), .ZN(net_187) );
INV_X4 inst_2079 ( .ZN(net_1628), .A(net_1626) );
OAI21_X4 inst_102 ( .ZN(net_2532), .A(net_2526), .B2(net_1640), .B1(net_982) );
DFFR_X2 inst_2527 ( .D(net_1642), .Q(net_1484), .CK(net_3061), .RN(x2480) );
INV_X2 inst_2231 ( .ZN(net_317), .A(net_316) );
CLKBUF_X2 inst_3277 ( .A(net_3234), .Z(net_3235) );
NAND2_X2 inst_1457 ( .ZN(net_1613), .A2(net_1612), .A1(net_1611) );
OAI21_X2 inst_144 ( .B2(net_1752), .ZN(net_1375), .A(net_1374), .B1(net_280) );
INV_X8 inst_1818 ( .A(net_2587), .ZN(net_2269) );
NAND2_X2 inst_1438 ( .A1(net_1687), .A2(net_1561), .ZN(net_1441) );
AOI21_X2 inst_2786 ( .B1(net_1363), .A(net_717), .ZN(net_438), .B2(net_394) );
NAND2_X2 inst_1224 ( .A1(net_1585), .A2(net_1532), .ZN(net_692) );
INV_X4 inst_1924 ( .A(net_848), .ZN(net_314) );
NAND2_X2 inst_1170 ( .ZN(net_105), .A1(net_86), .A2(x1014) );
INV_X8 inst_1766 ( .A(net_1248), .ZN(net_994) );
NAND2_X4 inst_880 ( .A2(net_2320), .ZN(net_1833), .A1(net_266) );
DFFR_X1 inst_2596 ( .D(net_2755), .CK(net_3418), .RN(x2480), .Q(x347) );
CLKBUF_X2 inst_2974 ( .A(net_2931), .Z(net_2932) );
CLKBUF_X2 inst_3022 ( .A(net_2952), .Z(net_2980) );
INV_X4 inst_1895 ( .ZN(net_426), .A(net_345) );
NAND3_X2 inst_680 ( .ZN(net_2510), .A3(net_2507), .A2(net_1287), .A1(net_1015) );
NAND2_X4 inst_785 ( .A2(net_2052), .ZN(net_1087), .A1(net_1081) );
AOI22_X2 inst_2730 ( .B1(net_2320), .ZN(net_1674), .A2(net_721), .B2(net_643), .A1(net_247) );
INV_X2 inst_2362 ( .ZN(net_1717), .A(net_1716) );
CLKBUF_X2 inst_3445 ( .A(net_3270), .Z(net_3403) );
CLKBUF_X2 inst_3299 ( .A(net_3256), .Z(net_3257) );
NAND2_X4 inst_737 ( .A1(net_2597), .ZN(net_613), .A2(net_234) );
CLKBUF_X2 inst_3255 ( .A(net_2944), .Z(net_3213) );
CLKBUF_X2 inst_2856 ( .A(net_2813), .Z(net_2814) );
NAND2_X4 inst_961 ( .ZN(net_2282), .A1(net_2280), .A2(net_848) );
NAND2_X4 inst_876 ( .A2(net_2269), .ZN(net_1790), .A1(net_1086) );
CLKBUF_X2 inst_2979 ( .A(net_2931), .Z(net_2937) );
NAND2_X2 inst_1590 ( .A2(net_2587), .ZN(net_2270), .A1(net_769) );
NAND4_X2 inst_545 ( .ZN(net_2142), .A1(net_2141), .A3(net_1372), .A4(net_1197), .A2(net_792) );
INV_X2 inst_2318 ( .A(net_873), .ZN(net_82) );
NOR2_X2 inst_399 ( .ZN(net_1043), .A2(net_1042), .A1(net_1041) );
NAND2_X2 inst_1388 ( .A2(net_1921), .ZN(net_1271), .A1(net_1268) );
NAND4_X2 inst_527 ( .A4(net_2576), .A2(net_2247), .ZN(net_1435), .A1(net_1207), .A3(net_1036) );
INV_X16 inst_2433 ( .ZN(net_2351), .A(net_2350) );
NOR2_X4 inst_226 ( .A2(net_1162), .ZN(net_905), .A1(net_904) );
AOI22_X4 inst_2699 ( .ZN(net_2674), .B2(net_2239), .A1(net_1942), .B1(net_243), .A2(net_242) );
NAND2_X2 inst_1180 ( .ZN(net_90), .A1(net_86), .A2(x793) );
NOR2_X2 inst_414 ( .A1(net_1286), .ZN(net_1225), .A2(net_532) );
DFFR_X2 inst_2480 ( .Q(net_1543), .D(net_333), .CK(net_3316), .RN(x2480) );
NAND4_X2 inst_531 ( .ZN(net_1901), .A2(net_1727), .A1(net_1726), .A4(net_1392), .A3(net_1257) );
NAND4_X1 inst_562 ( .A2(net_2531), .ZN(net_1792), .A3(net_1791), .A1(net_1309), .A4(net_294) );
AOI22_X2 inst_2737 ( .A2(net_2781), .ZN(net_2305), .A1(net_295), .B1(net_126), .B2(x2062) );
INV_X2 inst_2316 ( .A(net_1356), .ZN(net_852) );
NOR2_X4 inst_212 ( .A2(net_1814), .ZN(net_486), .A1(net_485) );
AOI22_X2 inst_2732 ( .A2(net_2758), .ZN(net_1966), .A1(net_295), .B1(net_126), .B2(x1262) );
NAND2_X2 inst_1299 ( .A2(net_2479), .A1(net_2478), .ZN(net_897) );
NAND4_X4 inst_499 ( .A4(net_1655), .ZN(net_1130), .A2(net_1129), .A1(net_1128), .A3(net_1127) );
CLKBUF_X2 inst_3396 ( .A(net_3011), .Z(net_3354) );
INV_X4 inst_1952 ( .A(net_2061), .ZN(net_607) );
NAND2_X2 inst_1372 ( .A2(net_1439), .ZN(net_1196), .A1(net_969) );
NAND2_X2 inst_1360 ( .A1(net_1151), .ZN(net_1147), .A2(net_1145) );
NAND3_X2 inst_674 ( .ZN(net_2343), .A3(net_2342), .A2(net_2341), .A1(net_2340) );
INV_X2 inst_2400 ( .ZN(net_2570), .A(net_2569) );
NAND2_X2 inst_1451 ( .A1(net_2287), .ZN(net_2050), .A2(net_800) );
NOR2_X2 inst_466 ( .ZN(net_2121), .A1(net_1178), .A2(net_1033) );
AOI21_X4 inst_2761 ( .B2(net_2138), .ZN(net_709), .B1(net_464), .A(net_385) );
NAND2_X4 inst_989 ( .ZN(net_2425), .A2(net_2424), .A1(net_2423) );
INV_X2 inst_2283 ( .ZN(net_44), .A(x876) );
INV_X2 inst_2253 ( .A(net_1564), .ZN(net_148) );
CLKBUF_X2 inst_3038 ( .A(net_2995), .Z(net_2996) );
CLKBUF_X2 inst_2966 ( .A(net_2923), .Z(net_2924) );
INV_X4 inst_2009 ( .ZN(net_1000), .A(net_999) );
CLKBUF_X2 inst_3246 ( .A(net_3203), .Z(net_3204) );
NAND2_X4 inst_858 ( .A1(net_2043), .ZN(net_1687), .A2(net_373) );
CLKBUF_X2 inst_2868 ( .A(net_2825), .Z(net_2826) );
NAND2_X2 inst_1109 ( .A2(net_574), .ZN(net_260), .A1(net_231) );
NAND4_X4 inst_501 ( .A1(net_2715), .A2(net_2600), .ZN(net_1604), .A4(net_1603), .A3(net_793) );
INV_X4 inst_2093 ( .A(net_2647), .ZN(net_1725) );
NAND2_X2 inst_1081 ( .A1(net_2022), .ZN(net_457), .A2(net_376) );
CLKBUF_X2 inst_3195 ( .A(net_2893), .Z(net_3153) );
CLKBUF_X2 inst_3037 ( .A(net_2955), .Z(net_2995) );
INV_X2 inst_2381 ( .A(net_2424), .ZN(net_2025) );
CLKBUF_X2 inst_2936 ( .A(net_2865), .Z(net_2894) );
INV_X1 inst_2468 ( .ZN(net_2226), .A(net_2225) );
OAI21_X4 inst_54 ( .B1(net_1585), .ZN(net_622), .A(net_590), .B2(net_29) );
CLKBUF_X2 inst_2905 ( .A(net_2811), .Z(net_2863) );
INV_X8 inst_1832 ( .ZN(net_2404), .A(net_2403) );
NAND3_X4 inst_570 ( .A1(net_2355), .ZN(net_1657), .A2(net_1656), .A3(net_1655) );
AOI21_X2 inst_2819 ( .ZN(net_2566), .B2(net_2565), .B1(net_2563), .A(net_2558) );
NAND2_X2 inst_1570 ( .A2(net_2270), .ZN(net_2161), .A1(net_2053) );
NAND3_X2 inst_640 ( .A2(net_2266), .ZN(net_1710), .A3(net_1709), .A1(net_1708) );
NAND2_X2 inst_1482 ( .A2(net_2023), .A1(net_2001), .ZN(net_1728) );
NAND2_X2 inst_1420 ( .A1(net_1602), .ZN(net_1366), .A2(net_234) );
NAND2_X2 inst_1314 ( .A1(net_1717), .ZN(net_952), .A2(net_948) );
NAND2_X2 inst_1612 ( .ZN(net_2412), .A2(net_2239), .A1(net_245) );
NAND2_X2 inst_1478 ( .A1(net_2201), .ZN(net_1712), .A2(net_1184) );
NAND2_X2 inst_1156 ( .A2(net_1495), .ZN(net_125), .A1(net_117) );
CLKBUF_X2 inst_3378 ( .A(net_3335), .Z(net_3336) );
NAND2_X2 inst_1114 ( .A1(net_2239), .A2(net_825), .ZN(net_239) );
NOR2_X2 inst_454 ( .A1(net_2177), .A2(net_2111), .ZN(net_1998) );
NAND2_X4 inst_942 ( .ZN(net_2177), .A2(net_2176), .A1(net_849) );
INV_X4 inst_1880 ( .ZN(net_454), .A(net_387) );
NAND2_X2 inst_1295 ( .A2(net_1120), .A1(net_1068), .ZN(net_888) );
NOR2_X4 inst_262 ( .A1(net_1841), .ZN(net_1455), .A2(net_1422) );
INV_X4 inst_1982 ( .A(net_1136), .ZN(net_823) );
INV_X4 inst_2089 ( .A(net_2561), .ZN(net_1698) );
NAND4_X4 inst_497 ( .A1(net_2670), .A3(net_2534), .A2(net_2051), .A4(net_1993), .ZN(net_557) );
INV_X4 inst_1849 ( .A(net_2575), .ZN(net_518) );
NAND2_X2 inst_1679 ( .ZN(net_2718), .A2(net_1109), .A1(net_1108) );
INV_X4 inst_1976 ( .ZN(net_789), .A(net_526) );
INV_X4 inst_2195 ( .ZN(net_2707), .A(net_1583) );
AOI22_X2 inst_2744 ( .ZN(net_2410), .B2(net_1777), .B1(net_1564), .A1(net_616), .A2(net_210) );
INV_X4 inst_2168 ( .A(net_2444), .ZN(net_2443) );
NAND2_X4 inst_1035 ( .ZN(net_2710), .A1(net_1585), .A2(net_1531) );
INV_X2 inst_2215 ( .ZN(net_391), .A(net_390) );
NAND2_X2 inst_1335 ( .A2(net_1904), .ZN(net_1003), .A1(net_489) );
CLKBUF_X2 inst_3077 ( .A(net_3034), .Z(net_3035) );
INV_X4 inst_1855 ( .A(net_1035), .ZN(net_533) );
NOR2_X2 inst_337 ( .A1(net_2514), .ZN(net_505), .A2(net_363) );
INV_X2 inst_2384 ( .ZN(net_2159), .A(net_1181) );
CLKBUF_X2 inst_3128 ( .A(net_3085), .Z(net_3086) );
INV_X4 inst_1883 ( .A(net_1790), .ZN(net_380) );
NAND2_X2 inst_1212 ( .A1(net_1585), .A2(net_1529), .ZN(net_624) );
NAND2_X2 inst_1078 ( .ZN(net_461), .A1(net_460), .A2(net_374) );
NAND3_X2 inst_670 ( .ZN(net_2251), .A2(net_2248), .A3(net_1672), .A1(net_931) );
DFFR_X2 inst_2517 ( .D(net_2317), .Q(net_1503), .CK(net_2932), .RN(x2480) );
NAND2_X2 inst_1423 ( .A2(net_1577), .ZN(net_1376), .A1(net_586) );
INV_X16 inst_2419 ( .A(net_2360), .ZN(net_1927) );
NAND2_X4 inst_1034 ( .ZN(net_2711), .A2(net_2710), .A1(net_88) );
NOR2_X2 inst_418 ( .A1(net_2296), .ZN(net_1336), .A2(net_384) );
NAND2_X4 inst_864 ( .ZN(net_1711), .A2(net_1185), .A1(net_754) );
NAND2_X2 inst_1207 ( .A2(net_1007), .A1(net_927), .ZN(net_610) );
OAI21_X4 inst_86 ( .B2(net_2509), .ZN(net_2081), .B1(net_2080), .A(net_2079) );
NAND2_X4 inst_949 ( .ZN(net_2202), .A2(net_2167), .A1(net_1216) );
CLKBUF_X2 inst_3283 ( .A(net_3240), .Z(net_3241) );
NAND3_X2 inst_613 ( .A3(net_2695), .A1(net_1547), .ZN(net_1238), .A2(net_1021) );
INV_X4 inst_1992 ( .A(net_1927), .ZN(net_861) );
NAND2_X4 inst_1039 ( .ZN(net_2724), .A2(net_1302), .A1(net_1301) );
NAND2_X4 inst_714 ( .A1(net_244), .ZN(net_211), .A2(net_210) );
INV_X2 inst_2396 ( .ZN(net_2447), .A(net_1058) );
CLKBUF_X2 inst_3005 ( .A(net_2961), .Z(net_2963) );
CLKBUF_X2 inst_2895 ( .A(net_2851), .Z(net_2853) );
NAND2_X2 inst_1428 ( .A2(net_2571), .ZN(net_1386), .A1(net_1385) );
NOR2_X2 inst_483 ( .ZN(net_2582), .A2(net_2581), .A1(net_2580) );
AOI22_X2 inst_2739 ( .ZN(net_2324), .B2(net_2323), .B1(net_2321), .A2(net_2320), .A1(net_2318) );
INV_X4 inst_2109 ( .ZN(net_1865), .A(net_1862) );
INV_X8 inst_1826 ( .ZN(net_2397), .A(net_2396) );
NOR2_X4 inst_259 ( .ZN(net_1430), .A2(net_1262), .A1(net_1261) );
NAND2_X2 inst_1046 ( .A1(net_2664), .A2(net_2661), .ZN(net_559) );
INV_X4 inst_2020 ( .A(net_1236), .ZN(net_1045) );
NOR2_X4 inst_246 ( .ZN(net_1193), .A2(net_1192), .A1(net_930) );
NAND2_X2 inst_1061 ( .A2(net_1904), .A1(net_1864), .ZN(net_512) );
NAND3_X2 inst_635 ( .ZN(net_1639), .A3(net_1638), .A2(net_981), .A1(net_391) );
NAND2_X2 inst_1177 ( .A1(net_98), .ZN(net_97), .A2(x730) );
AOI21_X2 inst_2820 ( .ZN(net_2632), .B1(net_2631), .B2(net_2455), .A(net_499) );
INV_X2 inst_2326 ( .ZN(net_983), .A(net_981) );
DFFR_X1 inst_2548 ( .QN(net_2796), .D(net_1749), .Q(net_1542), .CK(net_3353), .RN(x2480) );
NAND2_X4 inst_807 ( .A2(net_2433), .A1(net_2404), .ZN(net_1288) );
NAND2_X4 inst_705 ( .A1(net_1332), .ZN(net_514), .A2(net_415) );
INV_X2 inst_2404 ( .ZN(net_2636), .A(net_1595) );
OAI21_X4 inst_72 ( .B2(net_1976), .B1(net_1798), .ZN(net_1400), .A(net_842) );
NAND2_X4 inst_911 ( .A2(net_2514), .ZN(net_1995), .A1(net_1994) );
NAND2_X2 inst_1578 ( .ZN(net_2206), .A2(net_2204), .A1(net_2071) );
NAND4_X2 inst_519 ( .A4(net_2102), .ZN(net_1112), .A2(net_1089), .A3(net_594), .A1(net_593) );
NAND2_X2 inst_1666 ( .ZN(net_2688), .A2(net_608), .A1(net_413) );
NAND2_X2 inst_1634 ( .ZN(net_2542), .A1(net_2541), .A2(net_2529) );
NAND2_X4 inst_909 ( .ZN(net_1982), .A2(net_1981), .A1(net_1979) );
NAND2_X4 inst_1003 ( .ZN(net_2498), .A1(net_2497), .A2(net_866) );
DFFR_X2 inst_2484 ( .Q(net_1497), .D(net_698), .CK(net_3292), .RN(x2480) );
NAND2_X4 inst_735 ( .A1(net_1585), .A2(net_1507), .ZN(net_587) );
NAND2_X2 inst_1529 ( .A2(net_2629), .ZN(net_1976), .A1(net_1975) );
NAND2_X2 inst_1053 ( .A1(net_1871), .A2(net_850), .ZN(net_535) );
OAI21_X2 inst_115 ( .B2(net_1690), .ZN(net_257), .A(net_167), .B1(net_144) );
CLKBUF_X2 inst_2919 ( .A(net_2876), .Z(net_2877) );
NAND2_X2 inst_1653 ( .ZN(net_2613), .A2(net_951), .A1(net_949) );
NAND2_X4 inst_894 ( .ZN(net_1926), .A1(net_1802), .A2(net_1012) );
INV_X16 inst_2425 ( .A(net_2180), .ZN(net_2132) );
INV_X4 inst_1872 ( .A(net_467), .ZN(net_411) );
NAND2_X4 inst_994 ( .ZN(net_2462), .A1(net_2461), .A2(net_2399) );
AOI21_X4 inst_2774 ( .B1(net_2438), .ZN(net_1866), .B2(net_731), .A(net_366) );
CLKBUF_X2 inst_3045 ( .A(net_3002), .Z(net_3003) );
NOR2_X4 inst_239 ( .ZN(net_1133), .A2(net_1039), .A1(net_839) );
NAND2_X2 inst_1582 ( .A2(net_2295), .ZN(net_2217), .A1(net_384) );
INV_X4 inst_2080 ( .A(net_1962), .ZN(net_1632) );
INV_X4 inst_1879 ( .ZN(net_450), .A(net_387) );
NAND2_X2 inst_1193 ( .A2(net_2239), .ZN(net_579), .A1(net_185) );
CLKBUF_X2 inst_2984 ( .A(net_2941), .Z(net_2942) );
NAND2_X2 inst_1625 ( .ZN(net_2486), .A1(net_2481), .A2(net_1666) );
CLKBUF_X2 inst_3258 ( .A(net_3215), .Z(net_3216) );
INV_X4 inst_1863 ( .A(net_2022), .ZN(net_428) );
OAI21_X2 inst_175 ( .ZN(net_2576), .B2(net_2575), .B1(net_2574), .A(net_2570) );
NAND3_X2 inst_593 ( .A2(net_894), .A1(net_659), .ZN(net_596), .A3(net_578) );
INV_X2 inst_2223 ( .A(net_807), .ZN(net_362) );
INV_X4 inst_2135 ( .ZN(net_2140), .A(net_1294) );
INV_X8 inst_1737 ( .ZN(net_421), .A(net_384) );
CLKBUF_X2 inst_2995 ( .A(net_2952), .Z(net_2953) );
INV_X8 inst_1840 ( .ZN(net_2506), .A(net_2408) );
INV_X8 inst_1805 ( .A(net_2062), .ZN(net_2055) );
NAND3_X2 inst_601 ( .A1(net_1462), .A3(net_932), .ZN(net_883), .A2(net_612) );
OAI21_X2 inst_133 ( .B2(net_1998), .ZN(net_1059), .B1(net_1057), .A(net_365) );
NAND2_X2 inst_1263 ( .A2(net_2318), .A1(net_2133), .ZN(net_742) );
CLKBUF_X2 inst_3119 ( .A(net_3076), .Z(net_3077) );
NAND2_X4 inst_764 ( .A2(net_2538), .A1(net_1639), .ZN(net_920) );
INV_X8 inst_1773 ( .A(net_2165), .ZN(net_1181) );
NOR2_X2 inst_479 ( .ZN(net_2538), .A2(net_2523), .A1(net_716) );
AOI222_X1 inst_2752 ( .C1(net_736), .B1(net_721), .ZN(net_304), .C2(net_217), .A2(net_216), .B2(net_198), .A1(net_158) );
CLKBUF_X2 inst_3330 ( .A(net_3287), .Z(net_3288) );
INV_X2 inst_2344 ( .ZN(net_1373), .A(net_1371) );
NAND2_X2 inst_1547 ( .A1(net_2483), .ZN(net_2076), .A2(net_2068) );
OAI22_X2 inst_29 ( .A2(net_2801), .ZN(net_1622), .A1(net_169), .B1(net_156), .B2(net_49) );
CLKBUF_X2 inst_3326 ( .A(net_3283), .Z(net_3284) );
NAND2_X1 inst_1721 ( .A2(net_1930), .A1(net_1796), .ZN(net_1643) );
NAND2_X2 inst_1583 ( .ZN(net_2223), .A1(net_2222), .A2(net_872) );
NAND2_X2 inst_1149 ( .A1(net_631), .A2(net_180), .ZN(net_166) );
NAND2_X4 inst_771 ( .A2(net_2408), .ZN(net_995), .A1(net_994) );
NAND2_X2 inst_1445 ( .ZN(net_1559), .A2(net_1558), .A1(net_1557) );
NAND2_X2 inst_1281 ( .A1(net_1849), .A2(net_1625), .ZN(net_832) );
NAND2_X2 inst_1509 ( .A2(net_2561), .ZN(net_1852), .A1(net_1407) );
CLKBUF_X2 inst_3088 ( .A(net_3045), .Z(net_3046) );
INV_X2 inst_2369 ( .A(net_2319), .ZN(net_1777) );
INV_X4 inst_2152 ( .A(net_2405), .ZN(net_2336) );
NAND2_X2 inst_1274 ( .A1(net_1800), .ZN(net_790), .A2(net_545) );
OAI21_X2 inst_126 ( .B1(net_1585), .ZN(net_871), .A(net_870), .B2(net_54) );
NAND2_X2 inst_1512 ( .ZN(net_1876), .A1(net_1873), .A2(net_302) );
NAND2_X2 inst_1631 ( .ZN(net_2514), .A1(net_2512), .A2(net_1905) );
NAND4_X2 inst_538 ( .ZN(net_1880), .A2(net_1879), .A1(net_1418), .A4(net_1108), .A3(net_1106) );
AND2_X4 inst_2831 ( .ZN(net_1891), .A2(net_688), .A1(net_186) );
DFFR_X1 inst_2651 ( .D(net_1542), .CK(net_3160), .RN(x2480), .Q(x20) );
NAND2_X2 inst_1319 ( .ZN(net_966), .A2(net_965), .A1(net_964) );
NAND2_X2 inst_1300 ( .A2(net_1169), .ZN(net_898), .A1(net_446) );
NAND2_X2 inst_1140 ( .A2(net_1943), .A1(net_645), .ZN(net_189) );
OAI22_X2 inst_35 ( .ZN(net_2487), .A1(net_2486), .B1(net_2481), .A2(net_2071), .B2(net_1069) );
NAND2_X4 inst_948 ( .A1(net_2721), .A2(net_2397), .ZN(net_2197) );
NAND2_X2 inst_1086 ( .A2(net_2567), .A1(net_2564), .ZN(net_420) );
NOR2_X2 inst_358 ( .A1(net_1915), .A2(net_807), .ZN(net_370) );
OAI21_X4 inst_48 ( .B1(net_2259), .A(net_641), .ZN(net_198), .B2(net_50) );
DFFR_X1 inst_2643 ( .D(net_1463), .CK(net_3220), .RN(x2480), .Q(x106) );
INV_X2 inst_2246 ( .A(net_2655), .ZN(net_168) );
INV_X8 inst_1756 ( .A(net_1585), .ZN(net_634) );
INV_X2 inst_2279 ( .ZN(net_48), .A(x990) );
NAND2_X1 inst_1688 ( .A1(net_1361), .ZN(net_443), .A2(net_442) );
NOR2_X2 inst_443 ( .A2(net_2424), .A1(net_2153), .ZN(net_1714) );
INV_X2 inst_2299 ( .ZN(net_29), .A(x997) );
DFFR_X1 inst_2600 ( .Q(net_2773), .D(net_1127), .CK(net_2970), .RN(x2480) );
INV_X8 inst_1800 ( .A(net_1921), .ZN(net_1920) );
INV_X4 inst_2038 ( .ZN(net_1194), .A(net_1192) );
INV_X4 inst_2044 ( .ZN(net_1234), .A(net_1233) );
NAND3_X2 inst_655 ( .A3(net_2520), .ZN(net_1974), .A1(net_674), .A2(net_496) );
NOR2_X2 inst_448 ( .A1(net_2114), .ZN(net_1840), .A2(net_1354) );
INV_X2 inst_2274 ( .ZN(net_53), .A(x748) );
NAND2_X1 inst_1700 ( .A2(net_2328), .ZN(net_186), .A1(net_185) );
DFFR_X1 inst_2571 ( .D(net_2767), .CK(net_3202), .RN(x2480), .Q(x83) );
NAND2_X4 inst_914 ( .ZN(net_2011), .A1(net_2010), .A2(net_1071) );
NAND3_X2 inst_695 ( .A1(net_2700), .ZN(net_2698), .A3(net_1408), .A2(net_1391) );
INV_X4 inst_2002 ( .A(net_1323), .ZN(net_944) );
NAND2_X4 inst_730 ( .A1(net_1585), .A2(net_1498), .ZN(net_114) );
NAND2_X2 inst_1642 ( .A2(net_2587), .ZN(net_2577), .A1(net_1083) );
NOR2_X2 inst_384 ( .A1(net_2521), .ZN(net_1214), .A2(net_1169) );
NAND2_X2 inst_1252 ( .A2(net_2131), .ZN(net_724), .A1(net_721) );
NOR2_X4 inst_321 ( .ZN(net_2554), .A2(net_1893), .A1(net_1892) );
NAND2_X2 inst_1343 ( .ZN(net_1055), .A2(net_1027), .A1(net_497) );
NAND3_X2 inst_608 ( .A2(net_2179), .A1(net_2111), .A3(net_2016), .ZN(net_1077) );
NAND2_X4 inst_834 ( .A2(net_1869), .ZN(net_1554), .A1(net_815) );
CLKBUF_X2 inst_2920 ( .A(net_2877), .Z(net_2878) );
DFFR_X2 inst_2493 ( .Q(net_1483), .D(net_694), .CK(net_2864), .RN(x2480) );
NAND2_X4 inst_966 ( .ZN(net_2317), .A2(net_2316), .A1(net_2315) );
CLKBUF_X2 inst_3185 ( .A(net_3142), .Z(net_3143) );
CLKBUF_X2 inst_2961 ( .A(net_2918), .Z(net_2919) );
NAND2_X2 inst_1246 ( .A2(net_1310), .ZN(net_695), .A1(net_694) );
NAND4_X2 inst_511 ( .ZN(net_749), .A2(net_748), .A4(net_501), .A1(net_500), .A3(net_443) );
OAI221_X2 inst_41 ( .B1(net_2264), .A(net_676), .C1(net_601), .C2(net_321), .ZN(net_320), .B2(net_319) );
NOR3_X4 inst_199 ( .A3(net_2440), .A1(net_2284), .A2(net_2118), .ZN(net_1685) );
CLKBUF_X2 inst_3131 ( .A(net_3088), .Z(net_3089) );
INV_X2 inst_2209 ( .A(net_938), .ZN(net_445) );
AOI22_X2 inst_2722 ( .ZN(net_1126), .A1(net_139), .B1(net_133), .B2(net_70), .A2(x2080) );
DFFR_X2 inst_2506 ( .D(net_2651), .Q(net_1495), .CK(net_2822), .RN(x2480) );
DFFR_X1 inst_2645 ( .D(net_1518), .CK(net_3258), .RN(x2480), .Q(x177) );
INV_X4 inst_1989 ( .A(net_2334), .ZN(net_846) );
NAND2_X2 inst_1164 ( .A1(net_2259), .A2(net_1465), .ZN(net_113) );
CLKBUF_X2 inst_3112 ( .A(net_3013), .Z(net_3070) );
OAI21_X2 inst_152 ( .ZN(net_1631), .B2(net_1361), .A(net_718), .B1(net_502) );
NAND2_X2 inst_1238 ( .ZN(net_663), .A1(net_98), .A2(x883) );
INV_X4 inst_2171 ( .ZN(net_2463), .A(net_2462) );
INV_X4 inst_2029 ( .ZN(net_1142), .A(net_1140) );
NAND2_X2 inst_1152 ( .A1(net_1585), .ZN(net_135), .A2(net_69) );
NAND2_X2 inst_1242 ( .A1(net_1970), .A2(net_1255), .ZN(net_678) );
CLKBUF_X2 inst_3402 ( .A(net_3354), .Z(net_3360) );
NAND2_X2 inst_1400 ( .A2(net_2454), .A1(net_1909), .ZN(net_1305) );
NAND2_X4 inst_1011 ( .ZN(net_2553), .A2(net_1456), .A1(net_1455) );
NAND4_X2 inst_540 ( .ZN(net_1925), .A1(net_1924), .A2(net_1149), .A3(net_1134), .A4(net_1133) );
INV_X2 inst_2356 ( .A(net_1646), .ZN(net_1645) );
NOR2_X2 inst_404 ( .ZN(net_1116), .A2(net_774), .A1(net_773) );
NAND2_X4 inst_998 ( .ZN(net_2473), .A1(net_2470), .A2(net_2068) );
CLKBUF_X2 inst_3209 ( .A(net_3166), .Z(net_3167) );
CLKBUF_X2 inst_3160 ( .A(net_2928), .Z(net_3118) );
OAI21_X4 inst_89 ( .ZN(net_2122), .A(net_1287), .B2(net_1205), .B1(net_996) );
CLKBUF_X2 inst_2861 ( .A(net_2818), .Z(net_2819) );
NAND2_X2 inst_1520 ( .ZN(net_1941), .A1(net_1258), .A2(x585) );
NOR2_X2 inst_388 ( .ZN(net_924), .A1(net_137), .A2(net_46) );
OAI21_X4 inst_66 ( .B2(net_2221), .B1(net_1279), .A(net_1218), .ZN(net_1157) );
CLKBUF_X2 inst_3216 ( .A(net_3173), .Z(net_3174) );
NAND2_X2 inst_1535 ( .A2(net_2177), .A1(net_2113), .ZN(net_1999) );
OAI21_X1 inst_182 ( .B2(net_2503), .ZN(net_147), .A(net_146), .B1(net_27) );
NOR2_X4 inst_273 ( .A2(net_2566), .ZN(net_1727), .A1(net_1256) );
NAND2_X4 inst_788 ( .ZN(net_1099), .A2(net_1098), .A1(net_586) );
NOR2_X2 inst_489 ( .ZN(net_2738), .A1(net_2736), .A2(net_1113) );
NAND2_X4 inst_931 ( .ZN(net_2110), .A2(net_1930), .A1(net_1796) );
CLKBUF_X2 inst_3174 ( .A(net_3131), .Z(net_3132) );
INV_X4 inst_1965 ( .ZN(net_744), .A(net_302) );
OAI211_X2 inst_192 ( .ZN(net_2491), .A(net_2490), .C2(net_2481), .B(net_1665), .C1(net_1644) );
NAND2_X2 inst_1674 ( .ZN(net_2709), .A1(net_2708), .A2(net_1584) );
INV_X16 inst_2418 ( .A(net_2327), .ZN(net_1689) );
NOR2_X2 inst_366 ( .A1(net_1728), .ZN(net_656), .A2(net_345) );
AOI22_X2 inst_2715 ( .A2(net_2762), .ZN(net_810), .A1(net_284), .B1(net_126), .B2(x1785) );
NAND2_X2 inst_1579 ( .ZN(net_2210), .A2(net_1943), .A1(net_1602) );
NAND2_X2 inst_1411 ( .A1(net_1435), .ZN(net_1341), .A2(net_1274) );
OAI21_X2 inst_149 ( .ZN(net_1584), .B1(net_1583), .A(net_868), .B2(net_557) );
OAI211_X2 inst_193 ( .B(net_2603), .ZN(net_2522), .C2(net_2518), .C1(net_673), .A(net_355) );
OAI221_X2 inst_39 ( .C2(net_1690), .A(net_735), .ZN(net_323), .B2(net_319), .B1(net_172), .C1(net_153) );
NAND2_X2 inst_1415 ( .A2(net_2627), .A1(net_2417), .ZN(net_1349) );
DFFR_X1 inst_2627 ( .Q(net_2770), .D(net_757), .CK(net_3024), .RN(x2480) );
NAND2_X1 inst_1709 ( .A2(net_856), .ZN(net_727), .A1(net_721) );
INV_X16 inst_2413 ( .A(net_1115), .ZN(net_716) );
NAND2_X2 inst_1574 ( .A2(net_2739), .ZN(net_2183), .A1(net_980) );
CLKBUF_X2 inst_3285 ( .A(net_2939), .Z(net_3243) );
CLKBUF_X2 inst_3301 ( .A(net_3072), .Z(net_3259) );
INV_X2 inst_2320 ( .A(net_2473), .ZN(net_890) );
CLKBUF_X2 inst_3173 ( .A(net_2859), .Z(net_3131) );
OAI21_X2 inst_125 ( .A(net_2363), .B2(net_2362), .ZN(net_862), .B1(net_861) );
NOR2_X4 inst_228 ( .ZN(net_939), .A1(net_268), .A2(net_241) );
DFFR_X2 inst_2534 ( .QN(net_2803), .D(net_1512), .CK(net_3152), .RN(x2480) );
NOR2_X2 inst_486 ( .ZN(net_2630), .A2(net_2628), .A1(net_568) );
INV_X2 inst_2202 ( .ZN(net_515), .A(net_514) );
CLKBUF_X2 inst_3180 ( .A(net_3137), .Z(net_3138) );
NAND2_X4 inst_707 ( .ZN(net_464), .A1(net_463), .A2(net_383) );
NAND2_X4 inst_1025 ( .ZN(net_2652), .A1(net_2651), .A2(net_823) );
NAND2_X2 inst_1240 ( .A1(net_2408), .A2(net_1632), .ZN(net_673) );
CLKBUF_X2 inst_2987 ( .A(net_2944), .Z(net_2945) );
NOR2_X4 inst_244 ( .A1(net_2029), .ZN(net_1187), .A2(net_1186) );
NAND2_X2 inst_1636 ( .ZN(net_2555), .A2(net_1459), .A1(net_544) );
AOI21_X2 inst_2804 ( .ZN(net_1221), .B1(net_1220), .A(net_1219), .B2(net_1218) );
NOR2_X2 inst_430 ( .A1(net_1460), .ZN(net_1422), .A2(net_1421) );
NAND2_X2 inst_1521 ( .A1(net_2320), .ZN(net_1945), .A2(net_198) );
DFFR_X1 inst_2576 ( .D(net_2763), .CK(net_3420), .RN(x2480), .Q(x331) );
NAND4_X2 inst_515 ( .A3(net_2630), .A1(net_2082), .A2(net_1801), .ZN(net_976), .A4(net_843) );
CLKBUF_X2 inst_3079 ( .A(net_2955), .Z(net_3037) );
DFFR_X1 inst_2631 ( .Q(net_2766), .D(net_1136), .CK(net_2947), .RN(x2480) );
NAND2_X2 inst_1501 ( .A2(net_2320), .ZN(net_1829), .A1(net_1828) );
DFFR_X1 inst_2563 ( .QN(net_2798), .Q(net_1536), .D(net_559), .CK(net_2973), .RN(x2480) );
NAND2_X4 inst_772 ( .A2(net_1768), .ZN(net_999), .A1(net_367) );
NAND2_X2 inst_1306 ( .A1(net_2237), .A2(net_1076), .ZN(net_918) );
HA_X1 inst_2473 ( .B(net_941), .A(net_605), .S(net_85), .CO(net_84) );
CLKBUF_X2 inst_3212 ( .A(net_3169), .Z(net_3170) );
NAND2_X1 inst_1698 ( .A2(net_2237), .A1(net_1410), .ZN(net_207) );
DFFR_X1 inst_2565 ( .D(net_1375), .Q(net_78), .CK(net_3077), .RN(x2480) );
NAND2_X4 inst_944 ( .ZN(net_2181), .A1(net_1597), .A2(net_1249) );
NAND2_X2 inst_1407 ( .A2(net_2040), .ZN(net_1324), .A1(net_905) );
CLKBUF_X2 inst_2945 ( .A(net_2902), .Z(net_2903) );
DFFR_X1 inst_2636 ( .D(net_79), .CK(net_3321), .RN(x2480), .Q(x152) );
NAND2_X2 inst_1584 ( .ZN(net_2227), .A2(net_2224), .A1(net_1695) );
NAND3_X2 inst_642 ( .A2(net_2555), .A1(net_2554), .ZN(net_1776), .A3(net_1775) );
NOR2_X2 inst_459 ( .ZN(net_2072), .A2(net_2068), .A1(net_1644) );
CLKBUF_X2 inst_2993 ( .A(net_2950), .Z(net_2951) );
CLKBUF_X2 inst_2864 ( .A(net_2821), .Z(net_2822) );
NAND2_X4 inst_1018 ( .ZN(net_2589), .A1(net_589), .A2(net_102) );
NOR2_X2 inst_445 ( .ZN(net_1784), .A2(net_1288), .A1(net_454) );
OAI21_X4 inst_93 ( .ZN(net_2231), .A(net_2230), .B1(net_431), .B2(net_393) );
CLKBUF_X2 inst_2933 ( .A(net_2890), .Z(net_2891) );
NAND3_X1 inst_700 ( .A2(net_2562), .A3(net_1934), .ZN(net_397), .A1(net_369) );
CLKBUF_X2 inst_3393 ( .A(net_2834), .Z(net_3351) );
NOR2_X2 inst_367 ( .A2(net_2562), .ZN(net_680), .A1(net_679) );
NAND3_X2 inst_606 ( .A1(net_2599), .ZN(net_990), .A3(net_989), .A2(net_988) );
CLKBUF_X2 inst_2942 ( .A(net_2899), .Z(net_2900) );
NAND2_X4 inst_957 ( .ZN(net_2244), .A2(net_1000), .A1(net_998) );
NAND2_X4 inst_853 ( .ZN(net_1672), .A1(net_1671), .A2(net_1172) );
NAND2_X4 inst_979 ( .ZN(net_2374), .A1(net_2219), .A2(net_1611) );
AOI22_X2 inst_2713 ( .A2(net_2771), .B1(net_296), .A1(net_279), .ZN(net_276), .B2(x1844) );
OAI21_X2 inst_139 ( .B2(net_2132), .A(net_1379), .ZN(net_1224), .B1(net_1010) );
NAND2_X4 inst_1008 ( .ZN(net_2537), .A1(net_2523), .A2(net_716) );
CLKBUF_X2 inst_3409 ( .A(net_3366), .Z(net_3367) );
NAND3_X2 inst_657 ( .A3(net_2722), .ZN(net_2034), .A2(net_1670), .A1(net_1599) );
NAND4_X1 inst_559 ( .A3(net_2243), .A1(net_1890), .A2(net_1575), .ZN(net_882), .A4(net_308) );
NAND2_X2 inst_1675 ( .ZN(net_2712), .A1(net_2711), .A2(net_2328) );
INV_X4 inst_1871 ( .A(net_1085), .ZN(net_530) );
NAND3_X2 inst_584 ( .A2(net_2565), .A1(net_2130), .A3(net_1815), .ZN(net_479) );
CLKBUF_X2 inst_3433 ( .A(net_2855), .Z(net_3391) );
NAND2_X2 inst_1316 ( .A2(net_2585), .A1(net_1064), .ZN(net_954) );
INV_X2 inst_2296 ( .ZN(net_32), .A(x1742) );
INV_X4 inst_2098 ( .A(net_2552), .ZN(net_1775) );
NOR2_X2 inst_470 ( .A2(net_2567), .ZN(net_2230), .A1(net_807) );
INV_X4 inst_1921 ( .ZN(net_296), .A(net_284) );
INV_X2 inst_2300 ( .ZN(net_28), .A(x2017) );
NOR2_X2 inst_450 ( .A1(net_2517), .A2(net_2401), .ZN(net_1972) );
NAND4_X2 inst_520 ( .ZN(net_1118), .A4(net_1117), .A1(net_1116), .A3(net_199), .A2(net_177) );
NAND2_X4 inst_745 ( .ZN(net_699), .A1(net_698), .A2(net_232) );
OAI21_X2 inst_148 ( .B1(net_2475), .A(net_2071), .ZN(net_1425), .B2(net_1419) );
CLKBUF_X2 inst_3405 ( .A(net_2967), .Z(net_3363) );
NAND4_X2 inst_554 ( .ZN(net_2626), .A2(net_2625), .A1(net_1896), .A3(net_1867), .A4(net_540) );
INV_X8 inst_1752 ( .A(net_1585), .ZN(net_98) );
OAI211_X2 inst_191 ( .B(net_2398), .A(net_2395), .ZN(net_2303), .C2(net_2098), .C1(net_2097) );
NAND2_X2 inst_1187 ( .A2(net_1021), .A1(net_686), .ZN(net_571) );
NAND2_X2 inst_1063 ( .A1(net_983), .ZN(net_500), .A2(net_499) );
INV_X4 inst_2032 ( .ZN(net_1164), .A(net_1163) );
AOI22_X2 inst_2700 ( .A2(net_2776), .ZN(net_316), .A1(net_283), .B1(net_126), .B2(x1435) );
DFFR_X1 inst_2638 ( .D(net_76), .CK(net_3246), .RN(x2480), .Q(x166) );
INV_X4 inst_1917 ( .A(net_1943), .ZN(net_321) );
OAI21_X4 inst_80 ( .B2(net_2075), .ZN(net_1846), .B1(net_1461), .A(net_1459) );
INV_X4 inst_2026 ( .ZN(net_1121), .A(net_1120) );
CLKBUF_X2 inst_3252 ( .A(net_3209), .Z(net_3210) );
NAND2_X4 inst_836 ( .A2(net_2433), .A1(net_2405), .ZN(net_1567) );
NAND2_X2 inst_1556 ( .ZN(net_2113), .A2(net_2112), .A1(net_2111) );
CLKBUF_X2 inst_3235 ( .A(net_3192), .Z(net_3193) );
NOR2_X4 inst_241 ( .A2(net_1821), .ZN(net_1148), .A1(net_433) );
NAND2_X2 inst_1059 ( .A2(net_2165), .ZN(net_520), .A1(net_448) );
NAND2_X2 inst_1075 ( .A2(net_2558), .ZN(net_471), .A1(net_439) );
NAND2_X4 inst_862 ( .A1(net_1934), .ZN(net_1697), .A2(net_1407) );
AOI222_X1 inst_2758 ( .C1(net_1943), .ZN(net_1830), .C2(net_1828), .A2(net_736), .B2(net_227), .A1(net_203), .B1(net_158) );
NAND2_X2 inst_1167 ( .ZN(net_108), .A1(net_86), .A2(x857) );
NAND2_X2 inst_1116 ( .A1(net_1260), .ZN(net_230), .A2(net_187) );
INV_X4 inst_2087 ( .ZN(net_1690), .A(net_1689) );
INV_X2 inst_2257 ( .ZN(net_121), .A(net_86) );
INV_X8 inst_1764 ( .A(net_1611), .ZN(net_836) );
INV_X4 inst_2184 ( .ZN(net_2618), .A(net_2616) );
NAND2_X4 inst_892 ( .A1(net_2749), .A2(net_2153), .ZN(net_1879) );
NAND2_X2 inst_1104 ( .A1(net_697), .ZN(net_331), .A2(net_235) );
NAND2_X2 inst_1303 ( .A1(net_2312), .A2(net_1823), .ZN(net_910) );
NAND2_X2 inst_1623 ( .ZN(net_2484), .A2(net_2481), .A1(net_1738) );
NAND2_X2 inst_1132 ( .A2(net_2237), .A1(net_246), .ZN(net_201) );
NAND2_X2 inst_1159 ( .A1(net_2503), .ZN(net_146), .A2(net_93) );
INV_X2 inst_2355 ( .ZN(net_1635), .A(net_282) );
CLKBUF_X2 inst_3136 ( .A(net_3093), .Z(net_3094) );
NOR2_X2 inst_402 ( .A1(net_1837), .ZN(net_1088), .A2(net_658) );
NAND2_X4 inst_819 ( .A1(net_2059), .ZN(net_1399), .A2(net_1012) );
NAND2_X4 inst_968 ( .ZN(net_2321), .A2(net_745), .A1(net_675) );
CLKBUF_X2 inst_3320 ( .A(net_3277), .Z(net_3278) );
NAND2_X2 inst_1468 ( .A1(net_2429), .A2(net_2362), .ZN(net_1678) );
CLKBUF_X2 inst_3452 ( .A(net_3409), .Z(net_3410) );
NAND2_X2 inst_1516 ( .ZN(net_1884), .A2(net_799), .A1(net_528) );
INV_X8 inst_1803 ( .A(net_2657), .ZN(net_1977) );
NOR2_X4 inst_329 ( .ZN(net_2667), .A2(net_2454), .A1(net_2453) );
NOR2_X1 inst_494 ( .ZN(net_2074), .A2(net_2068), .A1(net_1665) );
NAND3_X4 inst_574 ( .ZN(net_2198), .A1(net_2197), .A3(net_1739), .A2(net_1251) );
NAND2_X4 inst_938 ( .A1(net_2612), .ZN(net_2136), .A2(net_1319) );
CLKBUF_X2 inst_3153 ( .A(net_3110), .Z(net_3111) );
AOI21_X2 inst_2814 ( .A(net_2569), .B1(net_2390), .ZN(net_2242), .B2(net_2206) );
NOR2_X2 inst_386 ( .A1(net_1072), .ZN(net_917), .A2(net_915) );
DFFR_X1 inst_2617 ( .Q(net_2752), .D(net_235), .CK(net_3304), .RN(x2480) );
INV_X2 inst_2347 ( .A(net_1429), .ZN(net_1428) );
NAND2_X2 inst_1229 ( .A1(net_1585), .A2(net_1480), .ZN(net_646) );
NAND2_X4 inst_936 ( .ZN(net_2131), .A2(net_637), .A1(net_91) );
NAND2_X2 inst_1288 ( .ZN(net_1897), .A1(net_1585), .A2(net_1488) );
CLKBUF_X2 inst_3068 ( .A(net_3025), .Z(net_3026) );
CLKBUF_X2 inst_2894 ( .A(net_2851), .Z(net_2852) );
INV_X2 inst_2358 ( .A(net_2726), .ZN(net_1650) );
INV_X4 inst_2125 ( .ZN(net_2008), .A(net_2007) );
AOI21_X4 inst_2778 ( .ZN(net_2253), .B1(net_2252), .B2(net_2028), .A(net_1104) );
INV_X2 inst_2277 ( .ZN(net_50), .A(x515) );
CLKBUF_X2 inst_2959 ( .A(net_2840), .Z(net_2917) );
NAND3_X2 inst_599 ( .ZN(net_878), .A3(net_877), .A2(net_876), .A1(net_874) );
NAND2_X4 inst_1033 ( .ZN(net_2714), .A2(net_2713), .A1(net_2712) );
NAND2_X2 inst_1683 ( .ZN(net_2740), .A1(net_2736), .A2(net_1115) );
CLKBUF_X2 inst_2962 ( .A(net_2869), .Z(net_2920) );
CLKBUF_X2 inst_3004 ( .A(net_2961), .Z(net_2962) );
NAND2_X2 inst_1348 ( .A2(net_2268), .ZN(net_1084), .A1(net_1083) );
DFFR_X1 inst_2647 ( .D(net_1472), .CK(net_3360), .RN(x2480), .Q(x208) );
INV_X4 inst_2102 ( .ZN(net_1806), .A(net_1804) );
INV_X8 inst_1748 ( .A(net_1008), .ZN(net_210) );
NAND4_X2 inst_541 ( .A4(net_2263), .ZN(net_1932), .A3(net_1024), .A1(net_912), .A2(net_610) );
NAND2_X4 inst_811 ( .A2(net_2726), .A1(net_1439), .ZN(net_1320) );
NOR3_X2 inst_208 ( .ZN(net_2208), .A1(net_2207), .A2(net_1029), .A3(net_1028) );
INV_X1 inst_2456 ( .A(net_2804), .ZN(net_605) );
NAND4_X4 inst_505 ( .A1(net_2532), .ZN(net_2143), .A2(net_1631), .A3(net_1569), .A4(net_828) );
NAND2_X2 inst_1365 ( .ZN(net_1165), .A2(net_768), .A1(net_485) );
AOI22_X2 inst_2710 ( .A2(net_2765), .ZN(net_280), .A1(net_279), .B1(net_278), .B2(x2167) );
CLKBUF_X2 inst_2887 ( .A(net_2844), .Z(net_2845) );
NAND2_X2 inst_1058 ( .A2(net_1820), .A1(net_1454), .ZN(net_521) );
NOR3_X4 inst_198 ( .ZN(net_1896), .A3(net_1395), .A2(net_1393), .A1(net_1016) );
INV_X4 inst_1869 ( .A(net_2297), .ZN(net_549) );
CLKBUF_X2 inst_3360 ( .A(net_3317), .Z(net_3318) );
NAND2_X4 inst_897 ( .A1(net_2317), .ZN(net_1936), .A2(net_766) );
NAND2_X2 inst_1371 ( .ZN(net_1190), .A2(net_86), .A1(x945) );
NAND2_X2 inst_1201 ( .A2(net_2326), .ZN(net_594), .A1(net_252) );
NAND2_X2 inst_1473 ( .A2(net_2323), .A1(net_1838), .ZN(net_1693) );
NAND2_X2 inst_1644 ( .ZN(net_2583), .A2(net_2086), .A1(net_1789) );
INV_X8 inst_1788 ( .A(net_2284), .ZN(net_1767) );
NAND2_X4 inst_784 ( .A2(net_2061), .ZN(net_1085), .A1(net_1083) );
NAND2_X2 inst_1272 ( .A2(net_1000), .ZN(net_783), .A1(net_509) );
CLKBUF_X2 inst_3237 ( .A(net_2882), .Z(net_3195) );
NAND3_X2 inst_632 ( .ZN(net_2452), .A2(net_1617), .A1(net_1616), .A3(net_1244) );
NAND3_X2 inst_636 ( .ZN(net_1659), .A3(net_1421), .A2(net_1200), .A1(net_836) );
NAND2_X2 inst_1264 ( .A1(net_2219), .A2(net_1611), .ZN(net_753) );
CLKBUF_X2 inst_2852 ( .A(x3333), .Z(net_2810) );
XOR2_X2 inst_0 ( .B(net_2418), .Z(net_129), .A(net_84) );
INV_X4 inst_1927 ( .ZN(net_237), .A(net_163) );
OAI211_X4 inst_184 ( .B(net_2437), .A(net_2436), .C1(net_1509), .ZN(net_982), .C2(net_981) );
INV_X8 inst_1847 ( .ZN(net_2739), .A(net_2736) );
CLKBUF_X2 inst_3461 ( .A(net_3390), .Z(net_3419) );
NAND3_X2 inst_690 ( .ZN(net_2660), .A3(net_2659), .A2(net_2658), .A1(net_1884) );
INV_X4 inst_1907 ( .ZN(net_302), .A(net_301) );
NOR2_X2 inst_433 ( .A2(net_2742), .ZN(net_1569), .A1(net_1568) );
INV_X4 inst_2025 ( .A(net_2165), .ZN(net_1110) );
INV_X4 inst_1983 ( .ZN(net_2015), .A(net_656) );
INV_X1 inst_2461 ( .ZN(net_1103), .A(net_1102) );
NAND2_X4 inst_732 ( .A1(net_2803), .ZN(net_569), .A2(x2269) );
INV_X4 inst_2178 ( .ZN(net_2524), .A(net_2523) );
INV_X4 inst_2192 ( .ZN(net_2686), .A(net_2685) );
NOR2_X4 inst_263 ( .A2(net_1598), .ZN(net_1456), .A1(net_1143) );
OAI211_X2 inst_185 ( .C2(net_1643), .ZN(net_528), .A(net_527), .C1(net_456), .B(net_410) );
INV_X4 inst_1948 ( .ZN(net_95), .A(x2242) );
INV_X4 inst_2114 ( .ZN(net_1918), .A(net_1813) );
OAI21_X4 inst_75 ( .ZN(net_2051), .B1(net_1995), .B2(net_459), .A(net_442) );
OAI21_X2 inst_166 ( .ZN(net_2254), .B1(net_1900), .B2(net_1454), .A(net_1232) );
AOI21_X2 inst_2784 ( .B1(net_860), .ZN(net_568), .B2(net_538), .A(net_532) );
OAI21_X4 inst_79 ( .ZN(net_1772), .A(net_1611), .B1(net_1030), .B2(net_890) );
OAI21_X4 inst_106 ( .ZN(net_2722), .B1(net_2721), .B2(net_2463), .A(net_2396) );
NOR2_X2 inst_422 ( .A1(net_2020), .A2(net_1579), .ZN(net_1357) );
DFFR_X1 inst_2583 ( .D(net_2774), .CK(net_3177), .RN(x2480), .Q(x10) );
INV_X2 inst_2243 ( .A(net_1688), .ZN(net_172) );
INV_X8 inst_1757 ( .ZN(net_679), .A(net_352) );
DFFR_X1 inst_2654 ( .D(net_1470), .CK(net_3155), .RN(x2480), .Q(x36) );
NAND2_X2 inst_1426 ( .A1(net_1793), .ZN(net_1382), .A2(net_293) );
NAND2_X2 inst_1475 ( .ZN(net_1706), .A2(net_1705), .A1(net_1704) );
CLKBUF_X2 inst_3090 ( .A(net_3047), .Z(net_3048) );
NAND2_X2 inst_1637 ( .ZN(net_2569), .A2(net_2219), .A1(net_836) );
NAND2_X2 inst_1352 ( .A2(net_2693), .A1(net_1181), .ZN(net_1104) );
NAND2_X2 inst_1605 ( .ZN(net_2366), .A2(net_2365), .A1(net_2364) );
INV_X2 inst_2261 ( .ZN(net_66), .A(x1835) );
CLKBUF_X2 inst_2975 ( .A(net_2914), .Z(net_2933) );
INV_X8 inst_1741 ( .A(net_2094), .ZN(net_341) );
NAND2_X4 inst_1024 ( .ZN(net_2647), .A2(net_2646), .A1(net_2033) );
INV_X2 inst_2232 ( .ZN(net_308), .A(net_307) );
CLKBUF_X2 inst_3390 ( .A(net_2810), .Z(net_3348) );
NAND2_X2 inst_1658 ( .ZN(net_2634), .A2(net_1052), .A1(net_901) );
CLKBUF_X2 inst_2930 ( .A(net_2887), .Z(net_2888) );
NAND2_X2 inst_1410 ( .A1(net_1341), .ZN(net_1339), .A2(net_1276) );
NAND2_X1 inst_1689 ( .A2(net_1650), .ZN(net_436), .A1(net_435) );
AND2_X2 inst_2846 ( .A1(net_2353), .ZN(net_1129), .A2(net_1097) );
CLKBUF_X2 inst_2859 ( .A(net_2816), .Z(net_2817) );
NOR2_X2 inst_397 ( .ZN(net_1020), .A1(net_878), .A2(net_306) );
NAND2_X2 inst_1448 ( .A2(net_2108), .ZN(net_1558), .A1(net_1554) );
NAND4_X4 inst_504 ( .A1(net_2324), .A3(net_2265), .ZN(net_1804), .A4(net_1621), .A2(net_1620) );
CLKBUF_X2 inst_3192 ( .A(net_3149), .Z(net_3150) );
INV_X8 inst_1733 ( .A(net_672), .ZN(net_387) );
NOR2_X2 inst_440 ( .A2(net_1905), .ZN(net_1640), .A1(net_1638) );
INV_X8 inst_1816 ( .ZN(net_2200), .A(net_2199) );
NAND2_X2 inst_1297 ( .A2(net_2323), .ZN(net_894), .A1(net_892) );
CLKBUF_X2 inst_3194 ( .A(net_3151), .Z(net_3152) );
INV_X32 inst_2199 ( .ZN(net_1008), .A(net_1007) );
NAND2_X4 inst_918 ( .ZN(net_2026), .A2(net_2025), .A1(net_2024) );
INV_X2 inst_2373 ( .A(net_1824), .ZN(net_1823) );
NAND2_X2 inst_1173 ( .ZN(net_103), .A1(net_86), .A2(x1031) );
CLKBUF_X2 inst_3381 ( .A(net_3338), .Z(net_3339) );
NAND2_X2 inst_1091 ( .A1(net_2695), .ZN(net_403), .A2(net_360) );
INV_X4 inst_1887 ( .A(net_2483), .ZN(net_361) );
CLKBUF_X2 inst_2908 ( .A(net_2865), .Z(net_2866) );
NAND2_X2 inst_1331 ( .A1(net_2711), .ZN(net_989), .A2(net_221) );
OAI21_X4 inst_52 ( .B1(net_1585), .ZN(net_619), .A(net_591), .B2(net_36) );
INV_X4 inst_2074 ( .ZN(net_1587), .A(net_1586) );
NAND2_X2 inst_1393 ( .A1(net_1766), .ZN(net_1292), .A2(net_1045) );
NAND3_X2 inst_668 ( .A2(net_2387), .ZN(net_2228), .A3(net_2006), .A1(net_1695) );
INV_X4 inst_1862 ( .A(net_508), .ZN(net_483) );
CLKBUF_X2 inst_3223 ( .A(net_3180), .Z(net_3181) );
NOR2_X4 inst_221 ( .ZN(net_697), .A1(net_274), .A2(net_254) );
NAND2_X2 inst_1236 ( .A1(net_1877), .ZN(net_660), .A2(net_586) );
CLKBUF_X2 inst_3049 ( .A(net_3006), .Z(net_3007) );
CLKBUF_X2 inst_3313 ( .A(net_3270), .Z(net_3271) );
NAND2_X2 inst_1672 ( .ZN(net_2697), .A2(net_701), .A1(net_554) );
CLKBUF_X2 inst_3349 ( .A(net_3306), .Z(net_3307) );
INV_X4 inst_2015 ( .ZN(net_1025), .A(net_1024) );
INV_X2 inst_2334 ( .A(net_2548), .ZN(net_1183) );
CLKBUF_X2 inst_3179 ( .A(net_2965), .Z(net_3137) );
INV_X16 inst_2429 ( .ZN(net_2239), .A(net_2236) );
DFFR_X1 inst_2545 ( .QN(net_2792), .Q(net_1472), .D(net_1339), .CK(net_3081), .RN(x2480) );
CLKBUF_X2 inst_3059 ( .A(net_3016), .Z(net_3017) );
CLKBUF_X2 inst_2970 ( .A(net_2927), .Z(net_2928) );
INV_X2 inst_2210 ( .A(net_2250), .ZN(net_429) );
AOI21_X4 inst_2768 ( .ZN(net_1298), .B1(net_1297), .A(net_1236), .B2(net_436) );
NAND2_X4 inst_754 ( .A1(net_2633), .ZN(net_772), .A2(net_499) );
INV_X8 inst_1835 ( .ZN(net_2440), .A(net_2119) );
CLKBUF_X2 inst_2937 ( .A(net_2894), .Z(net_2895) );
INV_X4 inst_1910 ( .ZN(net_269), .A(net_259) );
DFFR_X1 inst_2590 ( .Q(net_2776), .D(net_668), .CK(net_2994), .RN(x2480) );
CLKBUF_X2 inst_2913 ( .A(net_2837), .Z(net_2871) );
DFFR_X1 inst_2587 ( .D(net_2772), .CK(net_2898), .RN(x2480), .Q(x378) );
NAND3_X2 inst_687 ( .A1(net_2671), .ZN(net_2633), .A2(net_2631), .A3(net_771) );
INV_X2 inst_2319 ( .A(net_2035), .ZN(net_885) );
INV_X8 inst_1774 ( .ZN(net_1228), .A(net_1227) );
NAND3_X2 inst_621 ( .A2(net_2040), .ZN(net_1327), .A3(net_1326), .A1(net_905) );
CLKBUF_X2 inst_3295 ( .A(net_3252), .Z(net_3253) );
CLKBUF_X2 inst_3115 ( .A(net_3072), .Z(net_3073) );
DFFR_X1 inst_2560 ( .QN(net_2791), .Q(net_1470), .D(net_1349), .CK(net_2998), .RN(x2480) );
NAND2_X4 inst_985 ( .A1(net_2498), .ZN(net_2394), .A2(net_1760) );
CLKBUF_X2 inst_3219 ( .A(net_3176), .Z(net_3177) );
INV_X2 inst_2225 ( .A(net_1730), .ZN(net_369) );
NAND2_X4 inst_815 ( .A1(net_1913), .ZN(net_1359), .A2(net_340) );
CLKBUF_X2 inst_3031 ( .A(net_2844), .Z(net_2989) );
INV_X4 inst_2165 ( .A(net_2588), .ZN(net_2423) );
DFFR_X2 inst_2513 ( .D(net_2258), .Q(net_1525), .CK(net_2820), .RN(x2480) );
INV_X2 inst_2254 ( .A(net_616), .ZN(net_144) );
NAND2_X4 inst_875 ( .A1(net_2088), .ZN(net_1789), .A2(net_1764) );
NAND2_X2 inst_1257 ( .ZN(net_733), .A1(net_98), .A2(x1146) );
CLKBUF_X2 inst_3298 ( .A(net_3237), .Z(net_3256) );
CLKBUF_X2 inst_3081 ( .A(net_3038), .Z(net_3039) );
NAND2_X2 inst_1387 ( .ZN(net_1267), .A1(net_220), .A2(net_180) );
CLKBUF_X2 inst_2923 ( .A(net_2837), .Z(net_2881) );
INV_X4 inst_1991 ( .ZN(net_857), .A(net_856) );
AOI22_X2 inst_2707 ( .A2(net_2753), .ZN(net_301), .A1(net_284), .B1(net_278), .B2(x1681) );
INV_X4 inst_2069 ( .ZN(net_1555), .A(net_1554) );
INV_X2 inst_2365 ( .ZN(net_1741), .A(net_1278) );
NAND2_X2 inst_1117 ( .A1(net_2320), .A2(net_825), .ZN(net_228) );
INV_X4 inst_2108 ( .ZN(net_1848), .A(net_1847) );
CLKBUF_X2 inst_3066 ( .A(net_3023), .Z(net_3024) );
INV_X2 inst_2250 ( .ZN(net_229), .A(net_185) );
INV_X4 inst_2007 ( .ZN(net_975), .A(net_974) );
CLKBUF_X2 inst_2978 ( .A(net_2935), .Z(net_2936) );
AOI22_X2 inst_2725 ( .B2(net_2386), .ZN(net_1209), .A2(net_825), .A1(net_221), .B1(net_200) );
NOR2_X2 inst_413 ( .A2(net_1963), .ZN(net_1205), .A1(net_532) );
NOR2_X4 inst_334 ( .ZN(net_2748), .A2(net_2066), .A1(net_1872) );
NAND2_X2 inst_1610 ( .A1(net_2487), .ZN(net_2388), .A2(net_1619) );
INV_X4 inst_2187 ( .ZN(net_2648), .A(net_844) );
NAND2_X4 inst_859 ( .ZN(net_1688), .A1(net_113), .A2(net_89) );
NAND2_X4 inst_805 ( .A1(net_2506), .A2(net_2402), .ZN(net_1281) );
OAI22_X2 inst_25 ( .B2(net_2792), .ZN(net_813), .A1(net_156), .B1(net_126), .A2(net_47) );
CLKBUF_X2 inst_3323 ( .A(net_2834), .Z(net_3281) );
NOR2_X2 inst_354 ( .A1(net_1905), .A2(net_394), .ZN(net_390) );
INV_X4 inst_2019 ( .A(net_2374), .ZN(net_1040) );
NAND2_X2 inst_1145 ( .A2(net_1689), .A1(net_1191), .ZN(net_177) );
NAND2_X2 inst_1042 ( .A2(net_2146), .A1(net_2144), .ZN(net_563) );
DFFR_X2 inst_2500 ( .QN(net_2806), .D(net_1431), .CK(net_2938), .RN(x2480) );
OAI21_X4 inst_69 ( .B2(net_2198), .B1(net_1662), .ZN(net_1254), .A(net_810) );
NOR2_X2 inst_373 ( .A2(net_1318), .ZN(net_780), .A1(net_360) );
CLKBUF_X2 inst_3434 ( .A(net_3391), .Z(net_3392) );
CLKBUF_X2 inst_3056 ( .A(net_2956), .Z(net_3014) );
NAND2_X1 inst_1691 ( .A2(net_1351), .A1(net_715), .ZN(net_408) );
INV_X4 inst_1868 ( .A(net_1152), .ZN(net_503) );
NAND2_X4 inst_844 ( .ZN(net_1610), .A1(net_743), .A2(net_565) );
DFFR_X2 inst_2489 ( .Q(net_1500), .D(net_326), .CK(net_2870), .RN(x2480) );
NAND3_X2 inst_595 ( .A3(net_2514), .A2(net_1508), .ZN(net_755), .A1(net_671) );
DFFR_X1 inst_2609 ( .Q(net_2781), .D(net_1920), .CK(net_3035), .RN(x2480) );
OAI22_X2 inst_22 ( .B2(net_2783), .B1(net_1586), .ZN(net_235), .A1(net_137), .A2(net_34) );
DFFR_X1 inst_2556 ( .QN(net_2795), .Q(net_1534), .D(net_1198), .CK(net_3017), .RN(x2480) );
NAND2_X1 inst_1717 ( .A2(net_2505), .ZN(net_1177), .A1(net_387) );
INV_X2 inst_2340 ( .A(net_2404), .ZN(net_1283) );
NOR2_X2 inst_460 ( .ZN(net_2073), .A2(net_2068), .A1(net_1069) );
CLKBUF_X2 inst_3099 ( .A(net_3056), .Z(net_3057) );
NAND2_X2 inst_1455 ( .ZN(net_1605), .A2(net_667), .A1(net_666) );
CLKBUF_X2 inst_3204 ( .A(net_3161), .Z(net_3162) );
NAND2_X1 inst_1704 ( .A1(net_634), .ZN(net_106), .A2(x2183) );
DFFR_X2 inst_2497 ( .Q(net_1486), .D(net_711), .CK(net_2943), .RN(x2480) );
CLKBUF_X2 inst_2901 ( .A(net_2858), .Z(net_2859) );
NAND2_X4 inst_767 ( .A2(net_2726), .ZN(net_959), .A1(net_350) );
CLKBUF_X2 inst_3421 ( .A(net_3378), .Z(net_3379) );
OAI21_X2 inst_161 ( .ZN(net_2019), .A(net_2018), .B2(net_2017), .B1(net_1192) );
NAND4_X1 inst_560 ( .A2(net_1696), .A3(net_1099), .A1(net_1067), .ZN(net_919), .A4(net_918) );
CLKBUF_X2 inst_3356 ( .A(net_3237), .Z(net_3314) );
OAI22_X4 inst_16 ( .B2(net_2806), .B1(net_1589), .A1(net_1585), .ZN(net_618), .A2(net_68) );
NAND2_X4 inst_718 ( .A1(net_615), .ZN(net_246), .A2(net_90) );
AOI21_X2 inst_2808 ( .ZN(net_1371), .B1(net_1370), .B2(net_1323), .A(net_999) );
OAI21_X2 inst_156 ( .B1(net_2325), .ZN(net_1779), .A(net_575), .B2(net_140) );
NAND2_X4 inst_1029 ( .ZN(net_2687), .A1(net_2686), .A2(net_669) );
INV_X8 inst_1777 ( .A(net_1851), .ZN(net_1407) );
INV_X8 inst_1802 ( .ZN(net_1964), .A(net_1963) );
NAND2_X4 inst_950 ( .A1(net_2295), .ZN(net_2215), .A2(net_1824) );
NAND2_X2 inst_1068 ( .ZN(net_1919), .A1(net_956), .A2(net_606) );
NAND2_X4 inst_886 ( .ZN(net_1855), .A2(net_1193), .A1(net_345) );
CLKBUF_X2 inst_3442 ( .A(net_3399), .Z(net_3400) );
INV_X16 inst_2408 ( .A(net_2408), .ZN(net_343) );
CLKBUF_X2 inst_2982 ( .A(net_2939), .Z(net_2940) );
AOI22_X4 inst_2693 ( .B1(net_2321), .A2(net_2239), .A1(net_2131), .ZN(net_1778), .B2(net_1777) );
CLKBUF_X2 inst_3359 ( .A(net_3129), .Z(net_3317) );
NAND2_X2 inst_1218 ( .A1(net_1585), .A2(net_1538), .ZN(net_630) );
NAND2_X2 inst_1324 ( .ZN(net_972), .A2(net_969), .A1(net_944) );
NOR2_X2 inst_342 ( .A1(net_2392), .ZN(net_441), .A2(net_440) );
NAND4_X2 inst_526 ( .A1(net_2645), .A2(net_2643), .A4(net_1875), .ZN(net_1405), .A3(net_1404) );
INV_X4 inst_2147 ( .ZN(net_2280), .A(net_2279) );
NAND2_X2 inst_1178 ( .ZN(net_96), .A1(net_86), .A2(x1063) );
INV_X4 inst_2091 ( .ZN(net_1702), .A(net_1697) );
NOR2_X2 inst_463 ( .ZN(net_2085), .A2(net_2084), .A1(net_2083) );
OAI21_X4 inst_96 ( .A(net_2567), .B1(net_2373), .ZN(net_2302), .B2(net_2096) );
NAND2_X2 inst_1534 ( .A2(net_2516), .A1(net_2338), .ZN(net_1990) );
CLKBUF_X2 inst_3104 ( .A(net_3034), .Z(net_3062) );
CLKBUF_X2 inst_3020 ( .A(net_2977), .Z(net_2978) );
OAI21_X4 inst_101 ( .B1(net_2632), .ZN(net_2528), .B2(net_2527), .A(net_2525) );
NAND2_X2 inst_1549 ( .ZN(net_2078), .A2(net_2068), .A1(net_1738) );
NOR2_X4 inst_319 ( .ZN(net_2519), .A2(net_2518), .A1(net_937) );
NAND2_X2 inst_1450 ( .ZN(net_1580), .A2(net_1578), .A1(net_426) );
INV_X16 inst_2422 ( .ZN(net_2068), .A(net_2067) );
CLKBUF_X2 inst_3123 ( .A(net_3080), .Z(net_3081) );
NAND3_X2 inst_649 ( .A3(net_2134), .ZN(net_1928), .A1(net_687), .A2(net_581) );
INV_X4 inst_1969 ( .A(net_1025), .ZN(net_757) );
CLKBUF_X2 inst_2881 ( .A(net_2838), .Z(net_2839) );
NAND2_X4 inst_821 ( .A1(net_2415), .ZN(net_1406), .A2(net_813) );
INV_X4 inst_2158 ( .ZN(net_2380), .A(net_2379) );
NAND2_X1 inst_1711 ( .ZN(net_748), .A1(net_522), .A2(net_390) );
CLKBUF_X2 inst_3426 ( .A(net_3383), .Z(net_3384) );
DFFR_X1 inst_2597 ( .D(net_2758), .CK(net_3121), .RN(x2480), .Q(x44) );
NAND4_X4 inst_500 ( .A4(net_2804), .A3(net_2419), .ZN(net_1585), .A2(net_81), .A1(net_80) );
NAND2_X4 inst_980 ( .ZN(net_2381), .A2(net_2380), .A1(net_2378) );
NAND2_X2 inst_1592 ( .A2(net_2567), .A1(net_2395), .ZN(net_2273) );
INV_X8 inst_1770 ( .ZN(net_1115), .A(net_1113) );
NAND4_X4 inst_510 ( .ZN(net_2642), .A1(net_2641), .A3(net_2163), .A4(net_2158), .A2(net_2154) );
INV_X4 inst_2052 ( .A(net_2406), .ZN(net_1287) );
NAND4_X2 inst_550 ( .ZN(net_2434), .A1(net_2370), .A4(net_2368), .A2(net_2367), .A3(net_1861) );
NAND2_X4 inst_995 ( .ZN(net_2466), .A1(net_2465), .A2(net_1990) );
NAND2_X2 inst_1575 ( .ZN(net_2188), .A2(net_2187), .A1(net_511) );
CLKBUF_X2 inst_3413 ( .A(net_2873), .Z(net_3371) );
INV_X1 inst_2470 ( .ZN(net_2278), .A(net_2276) );
INV_X16 inst_2436 ( .ZN(net_2386), .A(net_2236) );
AND2_X4 inst_2832 ( .ZN(net_1892), .A1(net_1432), .A2(net_690) );
NAND2_X2 inst_1677 ( .ZN(net_2717), .A1(net_2716), .A2(net_276) );
NAND2_X2 inst_1258 ( .A1(net_2326), .A2(net_2030), .ZN(net_734) );
NAND3_X2 inst_603 ( .A3(net_1510), .ZN(net_950), .A2(net_861), .A1(net_805) );
NAND2_X4 inst_830 ( .A2(net_2360), .ZN(net_1453), .A1(net_1452) );
CLKBUF_X2 inst_3141 ( .A(net_3098), .Z(net_3099) );
INV_X8 inst_1785 ( .A(net_2726), .ZN(net_1648) );
NOR2_X4 inst_291 ( .ZN(net_2105), .A2(net_2104), .A1(net_2103) );
CLKBUF_X2 inst_2878 ( .A(net_2831), .Z(net_2836) );
INV_X4 inst_1957 ( .ZN(net_684), .A(net_82) );
CLKBUF_X2 inst_3150 ( .A(net_3107), .Z(net_3108) );
DFFR_X2 inst_2494 ( .D(net_2378), .Q(net_1466), .CK(net_3216), .RN(x2480) );
NAND2_X2 inst_1060 ( .ZN(net_2049), .A2(net_1046), .A1(net_483) );
NAND2_X4 inst_776 ( .A2(net_1988), .A1(net_1571), .ZN(net_1038) );
DFFR_X1 inst_2661 ( .D(net_869), .CK(net_3233), .RN(x2480), .Q(x90) );
NAND2_X4 inst_900 ( .ZN(net_1948), .A2(net_1947), .A1(net_1946) );
NAND2_X2 inst_1419 ( .A2(net_1912), .ZN(net_1364), .A1(net_340) );
DFFR_X2 inst_2526 ( .Q(net_1523), .D(net_1270), .CK(net_3313), .RN(x2480) );
INV_X2 inst_2286 ( .ZN(net_41), .A(x780) );
NAND2_X4 inst_866 ( .A2(net_2362), .A1(net_2351), .ZN(net_1716) );
INV_X4 inst_2137 ( .ZN(net_2156), .A(net_2155) );
DFFR_X2 inst_2501 ( .QN(net_2807), .Q(net_1469), .D(net_328), .CK(net_3212), .RN(x2480) );
NAND2_X2 inst_1439 ( .A1(net_2005), .ZN(net_1442), .A2(net_300) );
INV_X4 inst_1972 ( .A(net_1937), .ZN(net_766) );
NAND4_X2 inst_558 ( .ZN(net_2702), .A4(net_2701), .A1(net_2700), .A3(net_1408), .A2(net_1391) );
AOI21_X2 inst_2807 ( .B2(net_1653), .ZN(net_1315), .B1(net_1314), .A(net_1313) );
NAND3_X2 inst_594 ( .A2(net_2454), .ZN(net_671), .A3(net_394), .A1(net_363) );
CLKBUF_X2 inst_2983 ( .A(net_2940), .Z(net_2941) );
INV_X4 inst_2175 ( .ZN(net_2507), .A(net_2505) );
NOR2_X4 inst_248 ( .ZN(net_1223), .A1(net_1222), .A2(net_959) );
NAND2_X2 inst_1632 ( .ZN(net_2531), .A2(net_2525), .A1(net_555) );
NAND2_X2 inst_1613 ( .ZN(net_2413), .A1(net_2323), .A2(net_209) );
CLKBUF_X2 inst_3107 ( .A(net_3064), .Z(net_3065) );
NOR2_X2 inst_389 ( .A2(net_2325), .A1(net_1733), .ZN(net_926) );
INV_X4 inst_1919 ( .A(net_1010), .ZN(net_252) );
NAND2_X4 inst_925 ( .ZN(net_2058), .A2(net_2057), .A1(net_2056) );
INV_X2 inst_2378 ( .ZN(net_1911), .A(net_1909) );
INV_X4 inst_2193 ( .ZN(net_2695), .A(net_2694) );
AOI22_X2 inst_2712 ( .A2(net_2770), .B1(net_296), .A1(net_279), .ZN(net_277), .B2(x1750) );
NAND2_X2 inst_1120 ( .A1(net_618), .ZN(net_222), .A2(net_221) );
NAND2_X2 inst_1382 ( .A2(net_2482), .ZN(net_1243), .A1(net_1072) );
AOI21_X2 inst_2795 ( .B2(net_2192), .A(net_2153), .ZN(net_904), .B1(net_584) );
NAND2_X2 inst_1141 ( .A1(net_244), .ZN(net_188), .A2(net_187) );
INV_X8 inst_1807 ( .ZN(net_2067), .A(net_1062) );
DFFR_X2 inst_2488 ( .D(net_1802), .Q(net_1539), .CK(net_3111), .RN(x2480) );
NAND2_X4 inst_881 ( .ZN(net_1836), .A2(net_1835), .A1(net_1834) );
NAND2_X2 inst_1536 ( .A1(net_2177), .ZN(net_2000), .A2(net_1351) );
NAND2_X4 inst_932 ( .A2(net_2443), .ZN(net_2120), .A1(net_2118) );
CLKBUF_X2 inst_3184 ( .A(net_3128), .Z(net_3142) );
OAI21_X2 inst_180 ( .ZN(net_2672), .B1(net_2667), .B2(net_1361), .A(net_389) );
NAND2_X4 inst_913 ( .A1(net_2271), .ZN(net_2004), .A2(net_1707) );
INV_X4 inst_1960 ( .ZN(net_698), .A(net_697) );
NAND2_X4 inst_731 ( .A1(net_635), .ZN(net_92), .A2(x675) );
NAND2_X4 inst_947 ( .ZN(net_2196), .A1(net_2195), .A2(net_2108) );
NAND2_X2 inst_1225 ( .A1(net_1585), .A2(net_1474), .ZN(net_640) );
INV_X1 inst_2459 ( .A(net_712), .ZN(net_711) );
NOR2_X2 inst_363 ( .A2(net_2327), .ZN(net_165), .A1(net_164) );
NOR2_X4 inst_301 ( .ZN(net_2248), .A2(net_2111), .A1(net_1351) );
INV_X4 inst_2141 ( .ZN(net_2195), .A(net_2193) );
NOR2_X4 inst_247 ( .A2(net_2377), .A1(net_1614), .ZN(net_1207) );
NOR2_X2 inst_403 ( .A1(net_1984), .ZN(net_1090), .A2(net_607) );
NOR2_X4 inst_302 ( .ZN(net_2252), .A2(net_1919), .A1(net_530) );
NAND3_X2 inst_673 ( .ZN(net_2334), .A1(net_1581), .A3(net_934), .A2(net_426) );
CLKBUF_X2 inst_3446 ( .A(net_3403), .Z(net_3404) );
CLKBUF_X2 inst_3287 ( .A(net_3244), .Z(net_3245) );
AOI22_X2 inst_2728 ( .A1(net_1826), .ZN(net_1513), .B1(net_112), .B2(net_76), .A2(x1490) );
NOR2_X4 inst_211 ( .A1(net_1451), .ZN(net_1216), .A2(net_970) );
DFFR_X2 inst_2483 ( .Q(net_1538), .D(net_334), .CK(net_3113), .RN(x2480) );
NAND2_X2 inst_1151 ( .A2(net_2237), .A1(net_631), .ZN(net_161) );
NAND2_X2 inst_1588 ( .ZN(net_2265), .A1(net_2262), .A2(net_221) );
CLKBUF_X2 inst_3120 ( .A(net_2841), .Z(net_3078) );
CLKBUF_X2 inst_2956 ( .A(net_2913), .Z(net_2914) );
NAND2_X2 inst_1414 ( .A1(net_1922), .ZN(net_1344), .A2(net_1343) );
NAND4_X1 inst_561 ( .ZN(net_1636), .A4(net_1635), .A1(net_1266), .A2(net_770), .A3(net_543) );
NOR2_X2 inst_449 ( .ZN(net_1886), .A2(net_1885), .A1(net_1883) );
NOR2_X2 inst_412 ( .A1(net_2074), .ZN(net_1201), .A2(net_1200) );
DFFR_X1 inst_2650 ( .D(net_1534), .CK(net_2843), .RN(x2480), .Q(x389) );
DFFR_X2 inst_2516 ( .D(net_2213), .Q(net_1520), .CK(net_2979), .RN(x2480) );
DFFR_X2 inst_2505 ( .Q(net_1515), .D(net_595), .CK(net_2936), .RN(x2480) );
AOI21_X2 inst_2790 ( .B2(net_2493), .B1(net_1645), .ZN(net_602), .A(net_449) );
INV_X4 inst_2138 ( .A(net_2273), .ZN(net_2168) );
INV_X4 inst_2155 ( .A(net_2362), .ZN(net_2349) );
NAND2_X2 inst_1506 ( .ZN(net_1844), .A1(net_126), .A2(x1933) );
NAND2_X2 inst_1641 ( .ZN(net_2579), .A2(net_2578), .A1(net_2577) );
NOR2_X2 inst_464 ( .ZN(net_2098), .A2(net_1915), .A1(net_362) );
AOI22_X2 inst_2736 ( .B1(net_2323), .A2(net_2237), .ZN(net_2057), .A1(net_1838), .B2(net_1688) );
NOR2_X2 inst_341 ( .A1(net_2120), .A2(net_685), .ZN(net_451) );
CLKBUF_X2 inst_3189 ( .A(net_3053), .Z(net_3147) );
CLKBUF_X2 inst_3249 ( .A(net_2989), .Z(net_3207) );
CLKBUF_X2 inst_3163 ( .A(net_3120), .Z(net_3121) );
NOR3_X4 inst_196 ( .ZN(net_901), .A3(net_900), .A1(net_804), .A2(net_652) );
DFFR_X2 inst_2504 ( .D(net_2434), .Q(net_1521), .CK(net_2826), .RN(x2480) );
NAND2_X2 inst_1567 ( .ZN(net_2152), .A1(net_2064), .A2(net_703) );
CLKBUF_X2 inst_3451 ( .A(net_3408), .Z(net_3409) );
INV_X2 inst_2359 ( .ZN(net_1663), .A(net_377) );
INV_X16 inst_2417 ( .ZN(net_1589), .A(net_1585) );
INV_X2 inst_2309 ( .A(net_1318), .ZN(net_779) );
NAND3_X2 inst_684 ( .ZN(net_2563), .A3(net_2562), .A1(net_2559), .A2(net_704) );
CLKBUF_X2 inst_3374 ( .A(net_3331), .Z(net_3332) );
NAND2_X2 inst_1403 ( .A2(net_2611), .A1(net_2440), .ZN(net_1318) );
CLKBUF_X2 inst_3438 ( .A(net_3395), .Z(net_3396) );
CLKBUF_X2 inst_3177 ( .A(net_3134), .Z(net_3135) );
NAND2_X2 inst_1361 ( .A2(net_1925), .ZN(net_1150), .A1(net_1147) );
NOR2_X4 inst_298 ( .ZN(net_2203), .A2(net_2202), .A1(net_2100) );
CLKBUF_X2 inst_3401 ( .A(net_3358), .Z(net_3359) );
INV_X4 inst_2180 ( .ZN(net_2558), .A(net_2557) );
INV_X4 inst_1856 ( .A(net_2217), .ZN(net_517) );
DFFR_X1 inst_2603 ( .Q(net_2763), .D(net_1987), .CK(net_3094), .RN(x2480) );
OAI221_X2 inst_42 ( .ZN(net_1378), .B2(net_1377), .C1(net_321), .A(net_291), .B1(net_285), .C2(net_168) );
INV_X4 inst_2153 ( .ZN(net_2338), .A(net_2337) );
INV_X2 inst_2208 ( .A(net_937), .ZN(net_446) );
NAND3_X2 inst_588 ( .A3(net_573), .ZN(net_290), .A1(net_251), .A2(net_236) );
NAND2_X2 inst_1479 ( .A2(net_2424), .ZN(net_1713), .A1(net_469) );
NAND2_X2 inst_1138 ( .A1(net_2328), .A2(net_200), .ZN(net_191) );
NAND2_X2 inst_1241 ( .A1(net_1585), .A2(net_1493), .ZN(net_675) );
NAND2_X4 inst_1038 ( .ZN(net_2725), .A2(net_2724), .A1(net_1303) );
INV_X4 inst_2040 ( .A(net_2603), .ZN(net_1218) );
NOR2_X2 inst_437 ( .ZN(net_1618), .A2(net_1421), .A1(net_835) );
INV_X4 inst_2174 ( .ZN(net_2500), .A(net_940) );
NAND2_X4 inst_940 ( .A2(net_2285), .ZN(net_2167), .A1(net_2166) );
NAND2_X4 inst_1004 ( .ZN(net_2515), .A1(net_2512), .A2(net_2454) );
CLKBUF_X2 inst_3201 ( .A(net_3158), .Z(net_3159) );
OAI211_X2 inst_189 ( .C1(net_2473), .ZN(net_2246), .C2(net_2219), .B(net_1660), .A(net_1659) );
NAND2_X2 inst_1356 ( .ZN(net_1122), .A2(net_1120), .A1(net_177) );
NAND2_X1 inst_1706 ( .A1(net_2239), .A2(net_1564), .ZN(net_573) );
DFFR_X1 inst_2628 ( .Q(net_2750), .D(net_2102), .CK(net_2951), .RN(x2480) );
INV_X1 inst_2450 ( .A(net_778), .ZN(net_379) );
OR2_X2 inst_14 ( .A2(net_2739), .ZN(net_1508), .A1(net_1363) );
INV_X4 inst_2196 ( .ZN(net_2715), .A(net_2714) );
INV_X2 inst_2220 ( .ZN(net_440), .A(net_369) );
NAND2_X2 inst_1045 ( .A1(net_882), .A2(net_881), .ZN(net_560) );
AOI22_X2 inst_2743 ( .ZN(net_2370), .A2(net_2239), .B1(net_2131), .B2(net_1689), .A1(net_645) );
NOR2_X4 inst_252 ( .ZN(net_1309), .A2(net_1308), .A1(net_749) );
NAND2_X4 inst_865 ( .ZN(net_1715), .A2(net_1712), .A1(net_1711) );
OAI21_X4 inst_62 ( .B1(net_1585), .ZN(net_927), .A(net_131), .B2(net_35) );
INV_X2 inst_2325 ( .A(net_2425), .ZN(net_968) );
INV_X4 inst_2083 ( .A(net_1858), .ZN(net_1652) );
NAND2_X4 inst_956 ( .ZN(net_2245), .A1(net_2244), .A2(net_1001) );
NAND2_X2 inst_1470 ( .A2(net_2379), .ZN(net_1686), .A1(net_1430) );
CLKBUF_X2 inst_2860 ( .A(x3333), .Z(net_2818) );
NOR2_X4 inst_251 ( .ZN(net_1300), .A2(net_597), .A1(net_596) );
NAND2_X2 inst_1074 ( .A1(net_611), .ZN(net_473), .A2(net_472) );
NAND2_X4 inst_879 ( .A2(net_2562), .A1(net_1918), .ZN(net_1815) );
INV_X2 inst_2247 ( .ZN(net_233), .A(net_158) );
NAND2_X2 inst_1213 ( .A1(net_1585), .A2(net_1525), .ZN(net_625) );
NAND2_X2 inst_1524 ( .ZN(net_1950), .A1(net_736), .A2(net_216) );
NAND2_X2 inst_1552 ( .ZN(net_2097), .A2(net_2095), .A1(net_1700) );
CLKBUF_X2 inst_3072 ( .A(net_3029), .Z(net_3030) );
NOR2_X2 inst_484 ( .ZN(net_2595), .A2(net_2594), .A1(net_1776) );
INV_X1 inst_2452 ( .A(net_621), .ZN(net_153) );
OAI22_X2 inst_32 ( .B2(net_2790), .ZN(net_2224), .B1(net_225), .A1(net_112), .A2(net_57) );
NOR2_X2 inst_428 ( .A1(net_2297), .ZN(net_1414), .A2(net_1413) );
INV_X8 inst_1821 ( .ZN(net_2295), .A(net_2294) );
NAND2_X2 inst_1602 ( .ZN(net_2342), .A2(net_2021), .A1(net_408) );
CLKBUF_X2 inst_3418 ( .A(net_3312), .Z(net_3376) );
NAND2_X4 inst_969 ( .A1(net_2504), .ZN(net_2322), .A2(x2242) );
NAND3_X2 inst_629 ( .ZN(net_1571), .A3(net_1570), .A1(net_1037), .A2(net_205) );
CLKBUF_X2 inst_3334 ( .A(net_3291), .Z(net_3292) );
NOR2_X2 inst_407 ( .A1(net_2401), .ZN(net_1168), .A2(net_343) );
NAND2_X2 inst_1100 ( .A2(net_2112), .ZN(net_715), .A1(net_345) );
DFFR_X2 inst_2528 ( .Q(net_1498), .D(net_1065), .CK(net_3122), .RN(x2480) );
NAND2_X4 inst_791 ( .A2(net_2705), .ZN(net_1140), .A1(net_1139) );
NAND2_X2 inst_1208 ( .A1(net_1335), .A2(net_849), .ZN(net_612) );
INV_X4 inst_2021 ( .ZN(net_1063), .A(net_468) );
OAI21_X4 inst_97 ( .ZN(net_2318), .A(net_648), .B2(net_599), .B1(net_598) );
NAND3_X2 inst_616 ( .A1(net_2510), .A3(net_2468), .ZN(net_1284), .A2(net_1281) );
CLKBUF_X2 inst_3383 ( .A(net_3119), .Z(net_3341) );
NAND2_X4 inst_898 ( .ZN(net_1944), .A2(net_1943), .A1(net_1942) );
NAND2_X2 inst_1191 ( .A2(net_2239), .ZN(net_576), .A1(net_198) );
INV_X8 inst_1793 ( .A(net_2259), .ZN(net_1826) );
INV_X4 inst_1977 ( .A(net_1672), .ZN(net_795) );
NAND2_X4 inst_775 ( .A2(net_2506), .ZN(net_1032), .A1(net_994) );
NAND4_X2 inst_533 ( .A1(net_2346), .A2(net_2299), .ZN(net_1753), .A4(net_1624), .A3(net_1623) );
DFFR_X2 inst_2478 ( .D(net_2686), .Q(net_1540), .CK(net_2922), .RN(x2480) );
NAND3_X2 inst_620 ( .A2(net_2619), .ZN(net_1322), .A3(net_1321), .A1(net_1105) );
NAND3_X2 inst_652 ( .ZN(net_1955), .A2(net_1334), .A3(net_827), .A1(net_826) );
INV_X8 inst_1784 ( .ZN(net_1641), .A(net_1638) );
CLKBUF_X2 inst_3118 ( .A(net_3075), .Z(net_3076) );
AOI222_X1 inst_2751 ( .A2(net_1942), .B2(net_1260), .C2(net_736), .B1(net_721), .ZN(net_305), .C1(net_198), .A1(net_158) );
INV_X8 inst_1760 ( .ZN(net_704), .A(net_341) );
INV_X4 inst_1874 ( .A(net_1320), .ZN(net_463) );
INV_X2 inst_2343 ( .A(net_2553), .ZN(net_1367) );
INV_X2 inst_2291 ( .ZN(net_37), .A(x843) );
INV_X4 inst_2071 ( .ZN(net_1566), .A(net_1565) );
NAND3_X2 inst_677 ( .ZN(net_2428), .A3(net_2427), .A2(net_2356), .A1(net_1648) );
OAI21_X2 inst_130 ( .B1(net_1585), .ZN(net_1024), .A(net_1023), .B2(net_32) );
NAND2_X2 inst_1427 ( .ZN(net_1383), .A2(net_895), .A1(net_189) );
DFFR_X1 inst_2538 ( .QN(net_2784), .Q(net_1517), .D(net_1405), .CK(net_3375), .RN(x2480) );
NAND2_X2 inst_1566 ( .ZN(net_2154), .A2(net_2153), .A1(net_2152) );
INV_X4 inst_2022 ( .ZN(net_1082), .A(net_1081) );
CLKBUF_X2 inst_3132 ( .A(net_2948), .Z(net_3090) );
AOI21_X2 inst_2821 ( .ZN(net_2639), .B1(net_2615), .A(net_1595), .B2(net_364) );
NAND2_X2 inst_1409 ( .ZN(net_1334), .A1(net_200), .A2(net_158) );
NAND2_X2 inst_1095 ( .A1(net_2454), .A2(net_1909), .ZN(net_358) );
INV_X16 inst_2439 ( .ZN(net_2481), .A(net_2480) );
OAI21_X2 inst_176 ( .ZN(net_2620), .B1(net_2618), .A(net_1110), .B2(net_1090) );
AND2_X4 inst_2826 ( .A2(net_2110), .A1(net_2016), .ZN(net_1335) );
INV_X2 inst_2242 ( .A(net_619), .ZN(net_181) );
OAI21_X4 inst_87 ( .B2(net_2397), .ZN(net_2089), .A(net_889), .B1(net_841) );
CLKBUF_X2 inst_2996 ( .A(net_2953), .Z(net_2954) );
NAND2_X2 inst_1054 ( .A1(net_1286), .ZN(net_534), .A2(net_533) );
NAND2_X2 inst_1332 ( .A1(net_1718), .ZN(net_992), .A2(net_948) );
NAND2_X2 inst_1336 ( .A1(net_1332), .ZN(net_1005), .A2(net_1004) );
CLKBUF_X2 inst_2918 ( .A(net_2858), .Z(net_2876) );
INV_X8 inst_1841 ( .ZN(net_2516), .A(net_2404) );
NAND2_X4 inst_972 ( .ZN(net_2346), .A1(net_1552), .A2(net_421) );
NAND2_X2 inst_1665 ( .ZN(net_2678), .A2(net_2677), .A1(net_2675) );
CLKBUF_X2 inst_3345 ( .A(net_3064), .Z(net_3303) );
AOI22_X2 inst_2721 ( .ZN(net_1119), .B1(net_633), .A1(net_115), .A2(net_75), .B2(x1769) );
CLKBUF_X2 inst_3264 ( .A(net_2958), .Z(net_3222) );
NAND2_X2 inst_1671 ( .ZN(net_2699), .A1(net_2698), .A2(net_310) );
CLKBUF_X2 inst_3074 ( .A(net_2899), .Z(net_3032) );
NAND2_X4 inst_800 ( .ZN(net_1245), .A1(net_1242), .A2(net_1062) );
INV_X8 inst_1843 ( .ZN(net_2518), .A(net_2517) );
NAND2_X4 inst_780 ( .ZN(net_1061), .A1(net_1060), .A2(net_160) );
OR2_X2 inst_10 ( .A2(net_1904), .ZN(net_903), .A1(net_802) );
INV_X2 inst_2332 ( .ZN(net_1079), .A(net_1077) );
OR2_X4 inst_4 ( .A2(net_2787), .ZN(net_781), .A1(net_634) );
CLKBUF_X2 inst_2884 ( .A(net_2841), .Z(net_2842) );
NAND3_X2 inst_600 ( .A3(net_2243), .A1(net_1890), .A2(net_1575), .ZN(net_880) );
CLKBUF_X2 inst_3272 ( .A(net_3029), .Z(net_3230) );
NAND2_X2 inst_1194 ( .A2(net_2239), .A1(net_618), .ZN(net_580) );
INV_X2 inst_2310 ( .A(net_1155), .ZN(net_787) );
NAND2_X2 inst_1089 ( .A1(net_704), .ZN(net_406), .A2(net_405) );
NOR3_X2 inst_204 ( .ZN(net_1293), .A1(net_1273), .A2(net_896), .A3(net_309) );
OAI21_X4 inst_49 ( .B2(net_2808), .B1(net_634), .ZN(net_216), .A(net_105) );
INV_X8 inst_1767 ( .A(net_2680), .ZN(net_1021) );
INV_X2 inst_2219 ( .A(net_679), .ZN(net_437) );
INV_X4 inst_1866 ( .A(net_995), .ZN(net_495) );
NAND2_X2 inst_1550 ( .ZN(net_2079), .A1(net_938), .A2(net_495) );
NAND4_X2 inst_546 ( .ZN(net_2214), .A2(net_2212), .A3(net_1781), .A1(net_1780), .A4(net_330) );
NAND2_X2 inst_1284 ( .A1(net_1361), .ZN(net_838), .A2(net_444) );
INV_X1 inst_2465 ( .ZN(net_1807), .A(net_1806) );
INV_X2 inst_2361 ( .A(net_2128), .ZN(net_1700) );
INV_X4 inst_1878 ( .A(net_2537), .ZN(net_529) );
NAND2_X4 inst_910 ( .ZN(net_1979), .A2(net_1978), .A1(net_1977) );
NAND2_X2 inst_1290 ( .ZN(net_870), .A2(net_869), .A1(net_137) );
NAND2_X4 inst_704 ( .ZN(net_539), .A1(net_538), .A2(net_409) );
NAND3_X2 inst_693 ( .ZN(net_2689), .A2(net_2688), .A3(net_2422), .A1(net_2421) );
INV_X2 inst_2226 ( .A(net_1351), .ZN(net_349) );
NAND2_X4 inst_765 ( .A2(net_1167), .ZN(net_937), .A1(net_382) );
NAND2_X2 inst_1276 ( .A1(net_1254), .A2(net_1253), .ZN(net_812) );
NOR2_X4 inst_256 ( .A1(net_1511), .ZN(net_1395), .A2(net_1394) );
NAND3_X2 inst_694 ( .ZN(net_2690), .A3(net_2164), .A2(net_481), .A1(net_386) );
INV_X4 inst_2046 ( .ZN(net_1250), .A(net_95) );
INV_X4 inst_1902 ( .ZN(net_334), .A(net_329) );
DFFR_X2 inst_2498 ( .Q(net_1541), .D(net_919), .CK(net_2957), .RN(x2480) );
NAND2_X4 inst_937 ( .ZN(net_2138), .A2(net_2137), .A1(net_2135) );
CLKBUF_X2 inst_3154 ( .A(net_2907), .Z(net_3112) );
NAND2_X4 inst_908 ( .A1(net_2283), .A2(net_2203), .ZN(net_1968) );
NOR2_X2 inst_355 ( .A1(net_1654), .A2(net_836), .ZN(net_375) );
NOR2_X4 inst_218 ( .A2(net_2055), .A1(net_1086), .ZN(net_661) );
CLKBUF_X2 inst_3422 ( .A(net_3189), .Z(net_3380) );
CLKBUF_X2 inst_2971 ( .A(net_2928), .Z(net_2929) );
NAND2_X2 inst_1342 ( .ZN(net_1054), .A1(net_927), .A2(net_736) );
CLKBUF_X2 inst_2967 ( .A(net_2887), .Z(net_2925) );
DFFR_X2 inst_2531 ( .QN(net_2805), .D(net_129), .CK(net_3108), .RN(x2480) );
NAND2_X4 inst_787 ( .ZN(net_1098), .A2(net_663), .A1(net_662) );
NAND2_X4 inst_1014 ( .ZN(net_2581), .A2(net_2165), .A1(net_1158) );
INV_X4 inst_2078 ( .A(net_2344), .ZN(net_1624) );
INV_X8 inst_1747 ( .A(net_1008), .ZN(net_221) );
NAND2_X4 inst_825 ( .A2(net_2489), .ZN(net_1434), .A1(net_1432) );
NAND2_X2 inst_1347 ( .ZN(net_1075), .A2(net_86), .A1(x523) );
DFFR_X1 inst_2586 ( .D(net_2753), .CK(net_3350), .RN(x2480), .Q(x229) );
NAND4_X4 inst_509 ( .ZN(net_2615), .A1(net_2614), .A2(net_2546), .A3(net_1600), .A4(net_950) );
NAND2_X2 inst_1656 ( .ZN(net_2623), .A1(net_2622), .A2(net_706) );
NAND2_X2 inst_1680 ( .ZN(net_2731), .A2(net_2730), .A1(net_1607) );
NAND3_X1 inst_699 ( .A2(net_2588), .A1(net_2271), .A3(net_583), .ZN(net_481) );
INV_X4 inst_1881 ( .A(net_718), .ZN(net_499) );
NAND2_X2 inst_1462 ( .ZN(net_1626), .A1(net_551), .A2(net_547) );
DFFR_X1 inst_2622 ( .Q(net_2758), .D(net_1014), .CK(net_3221), .RN(x2480) );
NAND2_X2 inst_1626 ( .ZN(net_2490), .A2(net_2481), .A1(net_1071) );
OAI21_X2 inst_153 ( .B1(net_2393), .A(net_2168), .B2(net_2128), .ZN(net_1699) );
INV_X2 inst_2273 ( .ZN(net_54), .A(x1333) );
CLKBUF_X2 inst_3034 ( .A(net_2991), .Z(net_2992) );
INV_X4 inst_1892 ( .A(net_1725), .ZN(net_414) );
DFFR_X1 inst_2574 ( .D(net_2756), .CK(net_2857), .RN(x2480), .Q(x413) );
NOR2_X4 inst_295 ( .ZN(net_2151), .A2(net_1458), .A1(net_1457) );
NAND2_X4 inst_726 ( .A2(net_692), .A1(net_691), .ZN(net_243) );
NAND2_X2 inst_1459 ( .A1(net_2073), .ZN(net_1617), .A2(net_1615) );
INV_X2 inst_2229 ( .A(net_934), .ZN(net_493) );
INV_X4 inst_2003 ( .A(net_2215), .ZN(net_948) );
NOR3_X2 inst_209 ( .ZN(net_2669), .A1(net_2668), .A3(net_1509), .A2(net_529) );
NAND2_X4 inst_964 ( .A2(net_2548), .ZN(net_2293), .A1(net_1679) );
AOI21_X2 inst_2787 ( .B1(net_2502), .A(net_684), .ZN(net_94), .B2(net_93) );
NAND2_X2 inst_1087 ( .A2(net_2406), .A1(net_532), .ZN(net_416) );
NOR2_X4 inst_320 ( .ZN(net_2551), .A1(net_2547), .A2(net_2429) );
INV_X8 inst_1781 ( .ZN(net_1439), .A(net_1438) );
CLKBUF_X2 inst_3372 ( .A(net_3329), .Z(net_3330) );
NAND3_X2 inst_607 ( .A2(net_1696), .A3(net_1100), .ZN(net_1068), .A1(net_1067) );
AOI21_X4 inst_2769 ( .B2(net_1914), .ZN(net_1358), .A(net_1356), .B1(net_824) );
DFFR_X1 inst_2599 ( .Q(net_2779), .D(net_2676), .CK(net_3099), .RN(x2480) );
INV_X16 inst_2432 ( .ZN(net_2327), .A(net_2323) );
INV_X16 inst_2426 ( .ZN(net_2179), .A(net_2176) );
NAND2_X2 inst_1245 ( .A2(net_2320), .ZN(net_688), .A1(net_621) );
NAND2_X2 inst_1375 ( .A2(net_1963), .ZN(net_1204), .A1(net_434) );
INV_X2 inst_2313 ( .A(net_1934), .ZN(net_809) );
XOR2_X1 inst_1 ( .B(net_2803), .Z(net_1512), .A(net_82) );
INV_X4 inst_1891 ( .A(net_2739), .ZN(net_444) );
NAND2_X2 inst_1485 ( .ZN(net_1734), .A2(net_1731), .A1(net_736) );
CLKBUF_X2 inst_3001 ( .A(net_2958), .Z(net_2959) );
AOI21_X2 inst_2818 ( .ZN(net_2496), .B2(net_2386), .A(net_1761), .B1(net_173) );
CLKBUF_X2 inst_3215 ( .A(net_3125), .Z(net_3173) );
NOR2_X4 inst_235 ( .A1(net_2019), .ZN(net_1080), .A2(net_1079) );
CLKBUF_X2 inst_3063 ( .A(net_3020), .Z(net_3021) );
CLKBUF_X2 inst_3008 ( .A(net_2874), .Z(net_2966) );
CLKBUF_X2 inst_3198 ( .A(net_2837), .Z(net_3156) );
DFFR_X1 inst_2564 ( .D(net_1401), .Q(net_77), .CK(net_3336), .RN(x2480) );
NOR2_X4 inst_317 ( .ZN(net_2488), .A2(net_2481), .A1(net_2205) );
NAND2_X4 inst_750 ( .ZN(net_745), .A1(net_635), .A2(x1086) );
INV_X8 inst_1812 ( .ZN(net_2137), .A(net_2136) );
NAND2_X2 inst_1123 ( .A1(net_1688), .A2(net_1009), .ZN(net_215) );
NAND2_X2 inst_1082 ( .A2(net_867), .A1(net_608), .ZN(net_452) );
CLKBUF_X2 inst_2904 ( .A(net_2861), .Z(net_2862) );
NOR2_X4 inst_278 ( .A1(net_2055), .ZN(net_1850), .A2(net_1706) );
INV_X2 inst_2383 ( .ZN(net_2682), .A(net_1029) );
NAND2_X1 inst_1701 ( .A1(net_169), .ZN(net_150), .A2(x1381) );
NOR2_X2 inst_467 ( .A2(net_2693), .ZN(net_2150), .A1(net_958) );
INV_X4 inst_1995 ( .A(net_2802), .ZN(net_873) );
OAI21_X4 inst_105 ( .ZN(net_2597), .B1(net_121), .A(net_118), .B2(net_40) );
CLKBUF_X2 inst_3456 ( .A(net_3405), .Z(net_3414) );
CLKBUF_X2 inst_2963 ( .A(net_2920), .Z(net_2921) );
NAND2_X2 inst_1628 ( .ZN(net_2501), .A2(net_2500), .A1(net_2499) );
NAND2_X2 inst_1329 ( .A2(net_1907), .ZN(net_987), .A1(net_342) );
INV_X1 inst_2469 ( .ZN(net_2264), .A(net_2262) );
NAND2_X2 inst_1204 ( .A1(net_643), .ZN(net_603), .A2(net_221) );
INV_X4 inst_2161 ( .ZN(net_2402), .A(net_2401) );
NOR2_X4 inst_225 ( .A2(net_2055), .A1(net_1086), .ZN(net_867) );
NAND3_X2 inst_625 ( .A3(net_2624), .A1(net_1699), .ZN(net_1402), .A2(net_1165) );
CLKBUF_X2 inst_3367 ( .A(net_3324), .Z(net_3325) );
AND2_X4 inst_2835 ( .ZN(net_1924), .A2(net_1146), .A1(net_1135) );
NAND4_X4 inst_508 ( .ZN(net_2414), .A4(net_2413), .A3(net_2412), .A2(net_2411), .A1(net_2410) );
NAND3_X4 inst_568 ( .A1(net_1591), .ZN(net_1060), .A3(net_689), .A2(net_267) );
NAND4_X2 inst_523 ( .A3(net_1691), .ZN(net_1268), .A1(net_1267), .A2(net_665), .A4(net_582) );
NAND2_X2 inst_1483 ( .A2(net_2647), .A1(net_2557), .ZN(net_1730) );
AOI22_X2 inst_2731 ( .A2(net_2774), .ZN(net_1740), .A1(net_283), .B1(net_126), .B2(x1192) );
INV_X2 inst_2207 ( .A(net_956), .ZN(net_448) );
NAND2_X2 inst_1492 ( .ZN(net_1755), .A1(net_1593), .A2(net_1366) );
OAI21_X2 inst_181 ( .ZN(net_2676), .B1(net_1585), .A(net_1330), .B2(net_31) );
DFFR_X1 inst_2618 ( .D(net_2750), .CK(net_3168), .RN(x2480), .Q(x57) );
NAND2_X2 inst_1135 ( .A1(net_2320), .A2(net_2131), .ZN(net_196) );
NAND3_X2 inst_590 ( .ZN(net_274), .A3(net_191), .A2(net_162), .A1(net_161) );
DFFR_X1 inst_2553 ( .QN(net_2786), .D(net_2542), .Q(net_1467), .CK(net_3421), .RN(x2480) );
NAND2_X4 inst_713 ( .A2(net_1121), .ZN(net_337), .A1(net_318) );
CLKBUF_X2 inst_3127 ( .A(net_3012), .Z(net_3085) );
CLKBUF_X2 inst_3042 ( .A(net_2999), .Z(net_3000) );
CLKBUF_X2 inst_2867 ( .A(net_2824), .Z(net_2825) );
CLKBUF_X2 inst_3243 ( .A(net_3200), .Z(net_3201) );
NAND2_X1 inst_1729 ( .ZN(net_2421), .A2(net_1329), .A1(net_475) );
CLKBUF_X2 inst_2898 ( .A(net_2855), .Z(net_2856) );
NAND2_X2 inst_1105 ( .ZN(net_287), .A2(net_265), .A1(net_223) );
CLKBUF_X2 inst_3398 ( .A(net_3018), .Z(net_3356) );
AOI22_X2 inst_2746 ( .A2(net_2755), .ZN(net_2540), .A1(net_295), .B1(net_126), .B2(x1877) );
NOR2_X2 inst_477 ( .ZN(net_2533), .A2(net_2526), .A1(net_525) );
NAND2_X4 inst_981 ( .ZN(net_2378), .A1(net_1891), .A2(net_939) );
NAND2_X2 inst_1266 ( .A1(net_1433), .ZN(net_763), .A2(net_762) );
NAND2_X2 inst_1368 ( .A2(net_1863), .ZN(net_1175), .A1(net_503) );
NOR2_X2 inst_423 ( .A1(net_2740), .ZN(net_1360), .A2(net_1359) );
NAND2_X4 inst_835 ( .ZN(net_1563), .A1(net_86), .A2(x497) );
CLKBUF_X2 inst_3305 ( .A(net_2930), .Z(net_3263) );
INV_X4 inst_2094 ( .A(net_2209), .ZN(net_1726) );
INV_X4 inst_2088 ( .ZN(net_1695), .A(net_1694) );
CLKBUF_X2 inst_3082 ( .A(net_3039), .Z(net_3040) );
NOR2_X4 inst_330 ( .ZN(net_2673), .A2(net_1953), .A1(net_1952) );
CLKBUF_X2 inst_3208 ( .A(net_3165), .Z(net_3166) );
CLKBUF_X2 inst_3417 ( .A(net_3374), .Z(net_3375) );
NAND2_X2 inst_1112 ( .A2(net_1076), .ZN(net_253), .A1(net_163) );
OAI21_X2 inst_165 ( .ZN(net_2163), .B2(net_2162), .B1(net_2161), .A(net_2160) );
NAND2_X4 inst_710 ( .A2(net_2023), .A1(net_816), .ZN(net_467) );
NAND2_X2 inst_1379 ( .A1(net_2427), .ZN(net_1222), .A2(net_1021) );
NAND2_X4 inst_941 ( .ZN(net_2169), .A1(net_683), .A2(net_430) );
CLKBUF_X2 inst_3350 ( .A(net_3307), .Z(net_3308) );
NOR2_X4 inst_271 ( .A2(net_2291), .A1(net_2245), .ZN(net_1683) );
INV_X2 inst_2393 ( .A(net_2694), .ZN(net_2439) );
NAND2_X2 inst_1176 ( .ZN(net_99), .A1(net_86), .A2(x956) );
INV_X8 inst_1817 ( .A(net_2587), .ZN(net_2267) );
INV_X8 inst_1838 ( .ZN(net_2489), .A(net_2481) );
OAI21_X4 inst_71 ( .B2(net_2623), .A(net_2396), .B1(net_1550), .ZN(net_1392) );
OAI21_X4 inst_56 ( .B1(net_1585), .ZN(net_631), .A(net_630), .B2(net_55) );
NOR2_X4 inst_308 ( .ZN(net_2311), .A1(net_1336), .A2(net_422) );
NAND2_X2 inst_1546 ( .ZN(net_2070), .A2(net_2068), .A1(net_1610) );
NAND2_X2 inst_1230 ( .A1(net_1585), .A2(net_1528), .ZN(net_648) );
NOR2_X2 inst_455 ( .ZN(net_2013), .A1(net_2009), .A2(net_1666) );
NAND2_X2 inst_1454 ( .A1(net_2237), .ZN(net_1603), .A2(net_1602) );
CLKBUF_X2 inst_2871 ( .A(net_2828), .Z(net_2829) );
NAND2_X2 inst_1232 ( .A1(net_1585), .A2(net_1535), .ZN(net_650) );
NAND2_X1 inst_1694 ( .ZN(net_264), .A2(net_246), .A1(net_158) );
CLKBUF_X2 inst_3231 ( .A(net_3188), .Z(net_3189) );
CLKBUF_X2 inst_3147 ( .A(net_3104), .Z(net_3105) );
DFFR_X1 inst_2540 ( .D(net_2709), .Q(net_72), .CK(net_3070), .RN(x2480) );
NAND2_X2 inst_1064 ( .A1(net_708), .A2(net_685), .ZN(net_498) );
INV_X4 inst_1945 ( .A(net_1258), .ZN(net_115) );
DFFR_X1 inst_2657 ( .D(net_1476), .CK(net_3190), .RN(x2480), .Q(x78) );
DFFR_X1 inst_2605 ( .D(net_2762), .CK(net_3398), .RN(x2480), .Q(x273) );
NAND2_X4 inst_758 ( .A1(net_2296), .A2(net_1824), .ZN(net_803) );
NOR2_X2 inst_336 ( .A2(net_993), .A1(net_806), .ZN(net_542) );
CLKBUF_X2 inst_3024 ( .A(net_2981), .Z(net_2982) );
NAND3_X4 inst_583 ( .ZN(net_2657), .A3(net_2656), .A1(net_1833), .A2(net_1832) );
INV_X4 inst_2146 ( .ZN(net_2276), .A(net_2275) );
INV_X4 inst_1904 ( .A(net_913), .ZN(net_318) );
CLKBUF_X2 inst_3437 ( .A(net_3394), .Z(net_3395) );
AOI22_X2 inst_2703 ( .A2(net_2779), .ZN(net_558), .A1(net_284), .B1(net_278), .B2(x1826) );
NOR2_X2 inst_376 ( .A1(net_2311), .ZN(net_804), .A2(net_802) );
INV_X4 inst_1939 ( .A(net_1585), .ZN(net_139) );
INV_X4 inst_2065 ( .ZN(net_1457), .A(net_530) );
CLKBUF_X2 inst_3085 ( .A(net_3042), .Z(net_3043) );
INV_X2 inst_2251 ( .A(net_212), .ZN(net_154) );
CLKBUF_X2 inst_3268 ( .A(net_3225), .Z(net_3226) );
CLKBUF_X2 inst_2902 ( .A(net_2816), .Z(net_2860) );
OAI21_X2 inst_143 ( .A(net_1619), .ZN(net_1355), .B2(net_1242), .B1(net_1241) );
INV_X4 inst_1953 ( .A(net_1585), .ZN(net_632) );
CLKBUF_X2 inst_3016 ( .A(net_2951), .Z(net_2974) );
INV_X4 inst_1958 ( .ZN(net_693), .A(net_290) );
INV_X2 inst_2337 ( .ZN(net_1895), .A(net_1597) );
CLKBUF_X2 inst_3250 ( .A(net_3207), .Z(net_3208) );
CLKBUF_X2 inst_3240 ( .A(net_3197), .Z(net_3198) );
INV_X8 inst_1778 ( .A(net_2219), .ZN(net_1421) );
INV_X8 inst_1736 ( .ZN(net_367), .A(net_350) );
CLKBUF_X2 inst_2943 ( .A(net_2900), .Z(net_2901) );
INV_X4 inst_1899 ( .A(net_1935), .ZN(net_352) );
NAND2_X4 inst_1040 ( .ZN(net_2734), .A1(net_333), .A2(net_248) );
NAND2_X2 inst_1593 ( .A2(net_2395), .ZN(net_2274), .A1(net_371) );
DFFR_X1 inst_2569 ( .D(net_2759), .CK(net_3229), .RN(x2480), .Q(x98) );
NAND2_X4 inst_724 ( .A2(net_2733), .A1(net_2732), .ZN(net_200) );
CLKBUF_X2 inst_3100 ( .A(net_3057), .Z(net_3058) );
AOI22_X2 inst_2716 ( .A2(net_2780), .ZN(net_830), .A1(net_295), .B1(net_126), .B2(x1915) );
INV_X1 inst_2449 ( .A(net_991), .ZN(net_386) );
CLKBUF_X2 inst_3228 ( .A(net_3185), .Z(net_3186) );
OAI21_X2 inst_111 ( .B2(net_2288), .A(net_2286), .ZN(net_509), .B1(net_508) );
NAND2_X2 inst_1596 ( .ZN(net_2308), .A2(net_2178), .A1(net_407) );
NAND2_X4 inst_975 ( .ZN(net_2359), .A2(net_1677), .A1(net_1676) );
CLKBUF_X2 inst_3146 ( .A(net_2946), .Z(net_3104) );
INV_X4 inst_2124 ( .ZN(net_2002), .A(net_115) );
NAND2_X1 inst_1723 ( .A1(net_2055), .ZN(net_1707), .A2(net_1706) );
CLKBUF_X2 inst_3278 ( .A(net_3235), .Z(net_3236) );
CLKBUF_X2 inst_3191 ( .A(net_3148), .Z(net_3149) );
AOI21_X2 inst_2789 ( .B1(net_1064), .B2(net_769), .ZN(net_584), .A(net_419) );
INV_X2 inst_2289 ( .ZN(net_93), .A(x2269) );
INV_X4 inst_2056 ( .ZN(net_1310), .A(net_1127) );
INV_X4 inst_2116 ( .ZN(net_1929), .A(net_1928) );
NAND2_X2 inst_1431 ( .A2(net_2000), .ZN(net_1394), .A1(net_746) );
NAND2_X2 inst_1435 ( .A2(net_1823), .ZN(net_1415), .A1(net_1412) );
INV_X2 inst_2265 ( .ZN(net_62), .A(x535) );
NOR2_X4 inst_284 ( .A1(net_1996), .ZN(net_1993), .A2(net_1992) );
NAND2_X2 inst_1398 ( .ZN(net_1303), .A1(net_1300), .A2(net_1299) );
AND2_X4 inst_2825 ( .A2(net_2693), .A1(net_2165), .ZN(net_850) );
NAND2_X2 inst_1555 ( .ZN(net_2106), .A1(net_150), .A2(net_124) );
NAND2_X2 inst_1293 ( .A1(net_2491), .ZN(net_884), .A2(net_418) );
DFFR_X1 inst_2579 ( .D(net_2769), .CK(net_3370), .RN(x2480), .Q(x201) );
NOR2_X4 inst_280 ( .A2(net_2360), .ZN(net_1863), .A1(net_1862) );
AND2_X2 inst_2849 ( .A1(net_2655), .A2(net_2320), .ZN(net_1868) );
AOI22_X2 inst_2750 ( .ZN(net_2747), .B2(net_2237), .B1(net_647), .A1(net_245), .A2(net_158) );
INV_X8 inst_1804 ( .ZN(net_2017), .A(net_2016) );
INV_X16 inst_2440 ( .ZN(net_2483), .A(net_2481) );
NOR2_X2 inst_346 ( .A1(net_2363), .A2(net_1819), .ZN(net_417) );
NAND2_X2 inst_1467 ( .ZN(net_1669), .A1(net_1668), .A2(net_525) );
DFFR_X1 inst_2640 ( .D(net_77), .CK(net_3136), .RN(x2480), .Q(x484) );
CLKBUF_X2 inst_3157 ( .A(net_3114), .Z(net_3115) );
NAND2_X4 inst_978 ( .ZN(net_2371), .A2(net_1725), .A1(net_485) );
NAND2_X1 inst_1713 ( .A1(net_2000), .A2(net_934), .ZN(net_820) );
CLKBUF_X2 inst_2955 ( .A(net_2898), .Z(net_2913) );
INV_X4 inst_2183 ( .ZN(net_2614), .A(net_2613) );
CLKBUF_X2 inst_3327 ( .A(net_3284), .Z(net_3285) );
DFFR_X1 inst_2659 ( .D(net_1501), .CK(net_3186), .RN(x2480), .Q(x64) );
CLKBUF_X2 inst_3137 ( .A(net_2908), .Z(net_3095) );
INV_X4 inst_2134 ( .ZN(net_2108), .A(net_2107) );
INV_X8 inst_1744 ( .A(net_629), .ZN(net_255) );
AND2_X4 inst_2834 ( .ZN(net_1922), .A1(net_783), .A2(net_553) );
NAND2_X2 inst_1155 ( .A2(net_1500), .A1(net_598), .ZN(net_127) );
NAND2_X2 inst_1513 ( .ZN(net_1883), .A2(net_1882), .A1(net_1059) );
DFFR_X1 inst_2566 ( .QN(net_2783), .D(net_1637), .Q(net_1518), .CK(net_3013), .RN(x2480) );
NOR2_X1 inst_495 ( .ZN(net_2503), .A1(net_2501), .A2(net_684) );
NOR3_X2 inst_207 ( .ZN(net_1810), .A1(net_1809), .A3(net_1740), .A2(net_1278) );
NAND2_X2 inst_1051 ( .A2(net_1296), .A1(net_571), .ZN(net_537) );
NAND2_X4 inst_951 ( .ZN(net_2218), .A1(net_752), .A2(net_695) );
CLKBUF_X2 inst_3321 ( .A(net_3278), .Z(net_3279) );
INV_X4 inst_1864 ( .A(net_472), .ZN(net_427) );
NAND2_X2 inst_1545 ( .A2(net_2425), .ZN(net_2065), .A1(net_2064) );
CLKBUF_X2 inst_3338 ( .A(net_3295), .Z(net_3296) );
CLKBUF_X2 inst_3224 ( .A(net_2845), .Z(net_3182) );
NOR2_X4 inst_333 ( .ZN(net_2706), .A2(net_868), .A1(net_557) );
CLKBUF_X2 inst_3043 ( .A(net_3000), .Z(net_3001) );
NAND2_X4 inst_712 ( .A1(net_2214), .A2(net_1630), .ZN(net_338) );
NAND2_X2 inst_1215 ( .A1(net_1585), .A2(net_1466), .ZN(net_627) );
OAI21_X2 inst_131 ( .B1(net_1681), .ZN(net_1052), .B2(net_515), .A(net_364) );
NOR2_X2 inst_406 ( .A2(net_1768), .ZN(net_1155), .A1(net_1154) );
NOR2_X4 inst_328 ( .ZN(net_2641), .A2(net_2151), .A1(net_2150) );
CLKBUF_X2 inst_3111 ( .A(net_3068), .Z(net_3069) );
NAND2_X2 inst_1359 ( .A2(net_2557), .A1(net_2394), .ZN(net_1137) );
OAI21_X4 inst_47 ( .ZN(net_212), .B1(net_130), .A(net_125), .B2(net_53) );
INV_X4 inst_2035 ( .A(net_1863), .ZN(net_1174) );
CLKBUF_X2 inst_3188 ( .A(net_3145), .Z(net_3146) );
AOI21_X4 inst_2764 ( .ZN(net_1016), .B1(net_820), .B2(net_819), .A(net_817) );
CLKBUF_X2 inst_3129 ( .A(net_3032), .Z(net_3087) );
NAND2_X4 inst_818 ( .A1(net_1577), .ZN(net_1379), .A2(net_1009) );
INV_X4 inst_1984 ( .A(net_1357), .ZN(net_824) );
CLKBUF_X2 inst_2893 ( .A(net_2850), .Z(net_2851) );
NAND3_X4 inst_573 ( .ZN(net_1957), .A1(net_1956), .A2(net_726), .A3(net_184) );
OAI21_X4 inst_100 ( .ZN(net_2478), .B1(net_2477), .B2(net_1629), .A(net_277) );
NAND2_X4 inst_921 ( .ZN(net_2036), .A2(net_2035), .A1(net_2034) );
NAND2_X2 inst_1453 ( .A2(net_2418), .ZN(net_1596), .A1(net_873) );
NOR2_X4 inst_279 ( .ZN(net_1860), .A2(net_1200), .A1(net_1006) );
CLKBUF_X2 inst_3387 ( .A(net_3344), .Z(net_3345) );
CLKBUF_X2 inst_3274 ( .A(net_3231), .Z(net_3232) );
CLKBUF_X2 inst_3178 ( .A(net_3135), .Z(net_3136) );
CLKBUF_X2 inst_3007 ( .A(net_2964), .Z(net_2965) );
OAI21_X4 inst_81 ( .B1(net_2617), .ZN(net_1873), .B2(net_968), .A(net_475) );
AND2_X2 inst_2840 ( .A2(net_1011), .ZN(net_935), .A1(net_785) );
NAND4_X2 inst_525 ( .A3(net_2302), .A4(net_2301), .A2(net_2300), .ZN(net_1338), .A1(net_1206) );
AOI21_X4 inst_2781 ( .A(net_2569), .ZN(net_2472), .B2(net_2471), .B1(net_1860) );
NAND2_X4 inst_790 ( .ZN(net_1111), .A1(net_595), .A2(net_315) );
NOR2_X2 inst_434 ( .A2(net_2474), .A1(net_2452), .ZN(net_1575) );
CLKBUF_X2 inst_3455 ( .A(net_3412), .Z(net_3413) );
NAND2_X4 inst_1009 ( .ZN(net_2541), .A2(net_2540), .A1(net_2539) );
NAND2_X4 inst_1032 ( .ZN(net_2708), .A2(net_2707), .A1(net_2706) );
NAND2_X4 inst_906 ( .A1(net_2277), .ZN(net_1962), .A2(net_1211) );
NAND2_X2 inst_1206 ( .A2(net_2061), .ZN(net_609), .A1(net_380) );
CLKBUF_X2 inst_2954 ( .A(net_2911), .Z(net_2912) );
DFFR_X1 inst_2598 ( .Q(net_2756), .D(net_1588), .CK(net_2989), .RN(x2480) );
NAND2_X2 inst_1248 ( .A1(net_2423), .A2(net_1158), .ZN(net_703) );
INV_X2 inst_2402 ( .ZN(net_2580), .A(net_2579) );
NAND2_X2 inst_1392 ( .ZN(net_1290), .A1(net_685), .A2(net_360) );
INV_X4 inst_2197 ( .ZN(net_2744), .A(net_2743) );
DFFR_X1 inst_2616 ( .Q(net_2777), .D(net_1937), .CK(net_3031), .RN(x2480) );
NAND2_X4 inst_733 ( .A2(net_2239), .ZN(net_577), .A1(net_227) );
CLKBUF_X2 inst_3466 ( .A(net_3423), .Z(net_3424) );
INV_X4 inst_1959 ( .ZN(net_696), .A(net_694) );
DFFR_X1 inst_2582 ( .D(net_2752), .CK(net_3267), .RN(x2480), .Q(x170) );
NAND2_X2 inst_1476 ( .ZN(net_1705), .A1(net_1514), .A2(net_997) );
OAI21_X2 inst_142 ( .B1(net_2023), .A(net_1859), .B2(net_1672), .ZN(net_1353) );
INV_X2 inst_2249 ( .A(net_618), .ZN(net_155) );
OAI21_X4 inst_78 ( .B1(net_1812), .ZN(net_1747), .B2(net_1746), .A(net_1740) );
NAND2_X2 inst_1487 ( .A2(net_1792), .ZN(net_1736), .A1(net_1382) );
AOI21_X2 inst_2813 ( .ZN(net_2185), .B2(net_2183), .A(net_720), .B1(net_671) );
INV_X4 inst_2113 ( .A(net_2567), .ZN(net_1916) );
INV_X2 inst_2269 ( .ZN(net_58), .A(x629) );
OAI21_X2 inst_177 ( .ZN(net_2625), .B1(net_1856), .A(net_852), .B2(net_462) );
INV_X8 inst_1820 ( .ZN(net_2296), .A(net_2295) );
INV_X2 inst_2390 ( .ZN(net_2261), .A(x506) );
NAND2_X4 inst_783 ( .A1(net_2086), .A2(net_1789), .ZN(net_1081) );
INV_X8 inst_1780 ( .A(net_1665), .ZN(net_1432) );
OAI211_X4 inst_183 ( .A(net_2506), .B(net_1632), .C1(net_864), .ZN(net_674), .C2(net_398) );
NAND2_X2 inst_1436 ( .ZN(net_1440), .A2(net_1439), .A1(net_1021) );
INV_X4 inst_1933 ( .A(net_1008), .ZN(net_234) );
INV_X4 inst_2014 ( .ZN(net_1015), .A(net_450) );
NAND2_X4 inst_852 ( .A2(net_1920), .ZN(net_1667), .A1(net_1269) );
NAND2_X2 inst_1142 ( .A1(net_1877), .ZN(net_567), .A2(net_187) );
INV_X8 inst_1758 ( .A(net_686), .ZN(net_685) );
NAND3_X2 inst_615 ( .ZN(net_1261), .A1(net_1199), .A3(net_1092), .A2(net_577) );
INV_X2 inst_2271 ( .ZN(net_56), .A(x808) );
NAND2_X2 inst_1474 ( .A2(net_2128), .ZN(net_1701), .A1(net_414) );
INV_X4 inst_2045 ( .A(net_2482), .ZN(net_1242) );
AOI21_X1 inst_2822 ( .A(net_2217), .B2(net_1174), .B1(net_700), .ZN(net_546) );
INV_X1 inst_2467 ( .ZN(net_1983), .A(net_1977) );
INV_X4 inst_1920 ( .A(net_284), .ZN(net_278) );
INV_X4 inst_1848 ( .A(net_1175), .ZN(net_524) );
NAND2_X2 inst_1381 ( .A2(net_1619), .ZN(net_1244), .A1(net_1243) );
INV_X4 inst_2031 ( .ZN(net_1159), .A(net_1158) );
NAND3_X2 inst_643 ( .A2(net_2531), .ZN(net_1793), .A3(net_1791), .A1(net_1309) );
NAND2_X2 inst_1311 ( .A1(net_2804), .A2(net_2803), .ZN(net_940) );
NAND3_X2 inst_697 ( .ZN(net_2728), .A1(net_2727), .A3(net_2427), .A2(net_360) );
CLKBUF_X2 inst_3415 ( .A(net_3372), .Z(net_3373) );
NOR2_X2 inst_487 ( .ZN(net_2663), .A1(net_2662), .A2(net_1854) );
NAND2_X2 inst_1640 ( .ZN(net_2575), .A2(net_2492), .A1(net_840) );
CLKBUF_X2 inst_3234 ( .A(net_3191), .Z(net_3192) );
DFFR_X1 inst_2639 ( .D(net_70), .CK(net_3141), .RN(x2480), .Q(x444) );
INV_X4 inst_2133 ( .A(net_2567), .ZN(net_2099) );
INV_X4 inst_2163 ( .ZN(net_2419), .A(net_2418) );
DFFR_X2 inst_2509 ( .D(net_1902), .Q(net_1482), .CK(net_3206), .RN(x2480) );
NOR2_X2 inst_338 ( .A1(net_1855), .A2(net_1672), .ZN(net_474) );
INV_X16 inst_2412 ( .ZN(net_658), .A(net_585) );
DFFR_X1 inst_2542 ( .D(net_832), .Q(net_73), .CK(net_3069), .RN(x2480) );
CLKBUF_X2 inst_3091 ( .A(net_3048), .Z(net_3049) );
INV_X2 inst_2214 ( .A(net_488), .ZN(net_400) );
NOR2_X2 inst_417 ( .ZN(net_1304), .A2(net_720), .A1(net_525) );
NAND3_X2 inst_671 ( .ZN(net_2330), .A3(net_1373), .A2(net_788), .A1(net_787) );
INV_X4 inst_1861 ( .ZN(net_431), .A(net_430) );
INV_X4 inst_1997 ( .A(net_1062), .ZN(net_915) );
DFFS_X2 inst_2474 ( .Q(net_1492), .D(net_147), .QN(net_27), .CK(net_3179), .SN(x2480) );
NAND2_X4 inst_1017 ( .ZN(net_2586), .A1(net_1705), .A2(net_1704) );
NAND3_X4 inst_579 ( .ZN(net_2284), .A1(net_1842), .A3(net_1217), .A2(net_767) );
OAI22_X2 inst_21 ( .B2(net_2798), .ZN(net_670), .A1(net_137), .B1(net_126), .A2(net_64) );
DFFR_X2 inst_2495 ( .Q(net_1485), .D(net_325), .CK(net_2916), .RN(x2480) );
INV_X2 inst_2297 ( .ZN(net_31), .A(x1817) );
CLKBUF_X2 inst_3341 ( .A(net_3298), .Z(net_3299) );
NOR2_X4 inst_281 ( .A1(net_2335), .ZN(net_1867), .A2(net_1866) );
CLKBUF_X2 inst_3236 ( .A(net_3193), .Z(net_3194) );
NAND3_X2 inst_698 ( .ZN(net_2749), .A1(net_2748), .A2(net_2620), .A3(net_399) );
INV_X8 inst_1836 ( .ZN(net_2454), .A(net_1907) );
CLKBUF_X2 inst_3394 ( .A(net_3351), .Z(net_3352) );
INV_X4 inst_2004 ( .A(net_2061), .ZN(net_957) );
CLKBUF_X2 inst_3408 ( .A(net_3365), .Z(net_3366) );
INV_X2 inst_2311 ( .ZN(net_791), .A(net_790) );
OAI21_X4 inst_88 ( .A(net_2231), .ZN(net_2092), .B1(net_486), .B2(net_440) );
CLKBUF_X2 inst_2857 ( .A(net_2814), .Z(net_2815) );
NOR2_X4 inst_220 ( .A2(net_2071), .A1(net_753), .ZN(net_690) );
NAND2_X2 inst_1317 ( .A2(net_2061), .A1(net_1850), .ZN(net_956) );
NAND2_X2 inst_1585 ( .ZN(net_2249), .A2(net_2248), .A1(net_934) );
CLKBUF_X2 inst_2863 ( .A(net_2818), .Z(net_2821) );
DFFR_X2 inst_2508 ( .Q(net_1506), .D(net_1060), .CK(net_2912), .RN(x2480) );
INV_X4 inst_2170 ( .ZN(net_2459), .A(net_2458) );
NOR2_X2 inst_360 ( .A2(net_2427), .A1(net_1648), .ZN(net_339) );
CLKBUF_X2 inst_2941 ( .A(net_2850), .Z(net_2899) );
NAND2_X4 inst_773 ( .ZN(net_1018), .A1(net_1017), .A2(net_558) );
NOR2_X4 inst_245 ( .ZN(net_1189), .A1(net_1188), .A2(net_288) );
CLKBUF_X2 inst_2946 ( .A(net_2847), .Z(net_2904) );
INV_X4 inst_1873 ( .A(net_780), .ZN(net_460) );
NAND3_X2 inst_624 ( .A1(net_2550), .ZN(net_1390), .A2(net_1389), .A3(net_1176) );
NOR2_X4 inst_260 ( .A1(net_1548), .ZN(net_1450), .A2(net_1320) );
NAND2_X2 inst_1129 ( .A2(net_2237), .A1(net_621), .ZN(net_205) );
NAND2_X4 inst_837 ( .ZN(net_1577), .A1(net_1576), .A2(net_107) );
OAI21_X2 inst_147 ( .ZN(net_1423), .A(net_1421), .B2(net_1419), .B1(net_916) );
NAND2_X4 inst_744 ( .A2(net_1449), .ZN(net_694), .A1(net_693) );
NOR2_X4 inst_313 ( .ZN(net_2458), .A1(net_2127), .A2(net_260) );
CLKBUF_X2 inst_3211 ( .A(net_2961), .Z(net_3169) );
NAND2_X2 inst_1676 ( .ZN(net_2713), .A1(net_1009), .A2(net_647) );
NAND2_X4 inst_1041 ( .ZN(net_2736), .A2(net_2735), .A1(net_2734) );
CLKBUF_X2 inst_3114 ( .A(net_3071), .Z(net_3072) );
INV_X4 inst_2086 ( .A(net_1948), .ZN(net_1666) );
DFFR_X1 inst_2637 ( .D(net_73), .CK(net_2897), .RN(x2480), .Q(x370) );
NOR2_X4 inst_236 ( .ZN(net_1089), .A1(net_1088), .A2(net_218) );
NAND4_X2 inst_553 ( .ZN(net_2606), .A3(net_2604), .A2(net_1922), .A1(net_1293), .A4(net_1292) );
OAI21_X4 inst_65 ( .B1(net_1562), .ZN(net_1141), .B2(net_1140), .A(net_299) );
CLKBUF_X2 inst_3331 ( .A(net_3288), .Z(net_3289) );
NAND4_X2 inst_536 ( .ZN(net_1812), .A1(net_1811), .A4(net_1743), .A3(net_1742), .A2(net_1741) );
CLKBUF_X2 inst_3172 ( .A(net_3129), .Z(net_3130) );
NAND2_X4 inst_986 ( .ZN(net_2401), .A1(net_1429), .A2(net_906) );
NOR2_X4 inst_242 ( .A2(net_2123), .ZN(net_1149), .A1(net_834) );
INV_X2 inst_2386 ( .ZN(net_2178), .A(net_2176) );
NAND2_X2 inst_1422 ( .A2(net_2595), .ZN(net_1368), .A1(net_1367) );
NAND4_X2 inst_516 ( .A3(net_2744), .A4(net_2591), .ZN(net_1013), .A1(net_935), .A2(net_784) );
INV_X2 inst_2258 ( .A(net_632), .ZN(net_112) );
OAI211_X2 inst_190 ( .ZN(net_2683), .A(net_2050), .B(net_2049), .C2(net_1767), .C1(net_510) );
NAND2_X2 inst_1186 ( .A1(net_635), .ZN(net_87), .A2(x543) );
NAND2_X2 inst_1267 ( .A1(net_1241), .A2(net_1040), .ZN(net_762) );
NAND2_X2 inst_1507 ( .ZN(net_1847), .A2(net_1846), .A1(net_1773) );
NAND2_X2 inst_1221 ( .A1(net_1585), .A2(net_1486), .ZN(net_654) );
NAND2_X1 inst_1727 ( .A1(net_2196), .A2(net_2194), .ZN(net_2109) );
INV_X8 inst_1753 ( .A(net_569), .ZN(net_80) );
INV_X4 inst_2027 ( .ZN(net_1120), .A(net_1119) );
CLKBUF_X2 inst_2926 ( .A(net_2883), .Z(net_2884) );
NAND2_X2 inst_1166 ( .A1(net_2259), .A2(net_1539), .ZN(net_110) );
OAI21_X2 inst_116 ( .ZN(net_179), .A(net_123), .B1(net_115), .B2(net_63) );
INV_X8 inst_1739 ( .A(net_2111), .ZN(net_655) );
NOR2_X2 inst_416 ( .A2(net_2427), .ZN(net_1264), .A1(net_1263) );
NAND2_X2 inst_1133 ( .A2(net_2320), .A1(net_631), .ZN(net_199) );
NAND2_X2 inst_1158 ( .ZN(net_123), .A1(net_115), .A2(net_79) );
NOR2_X2 inst_471 ( .ZN(net_2243), .A1(net_2242), .A2(net_763) );
INV_X4 inst_1870 ( .A(net_1720), .ZN(net_415) );
INV_X4 inst_2062 ( .ZN(net_1413), .A(net_1412) );
INV_X2 inst_2350 ( .A(net_2219), .ZN(net_1459) );
INV_X4 inst_2103 ( .ZN(net_1811), .A(net_1809) );
NAND2_X2 inst_1406 ( .ZN(net_1325), .A1(net_1324), .A2(net_297) );
CLKBUF_X2 inst_3404 ( .A(net_3361), .Z(net_3362) );
NAND4_X2 inst_542 ( .ZN(net_1989), .A4(net_1987), .A1(net_1570), .A2(net_1037), .A3(net_205) );
OAI21_X2 inst_128 ( .B2(net_1440), .A(net_971), .ZN(net_896), .B1(net_685) );
NAND2_X4 inst_896 ( .ZN(net_1931), .A1(net_1642), .A2(net_1025) );
NOR2_X2 inst_339 ( .A2(net_1567), .ZN(net_465), .A1(net_396) );
NOR2_X2 inst_351 ( .A2(net_2219), .A1(net_835), .ZN(net_418) );
INV_X16 inst_2445 ( .ZN(net_2727), .A(net_2726) );
DFFR_X1 inst_2608 ( .Q(net_2774), .D(net_848), .CK(net_3327), .RN(x2480) );
CLKBUF_X2 inst_3039 ( .A(net_2996), .Z(net_2997) );
NAND2_X4 inst_973 ( .ZN(net_2350), .A1(net_1960), .A2(net_1881) );
CLKBUF_X2 inst_3435 ( .A(net_3392), .Z(net_3393) );
CLKBUF_X2 inst_3058 ( .A(net_3015), .Z(net_3016) );
DFFR_X1 inst_2557 ( .D(net_561), .Q(net_70), .CK(net_3058), .RN(x2480) );
NOR2_X2 inst_461 ( .A1(net_2484), .ZN(net_2075), .A2(net_2068) );
CLKBUF_X2 inst_3218 ( .A(net_3175), .Z(net_3176) );
DFFR_X2 inst_2521 ( .QN(net_2808), .D(net_759), .CK(net_2929), .RN(x2480) );
NAND2_X4 inst_829 ( .ZN(net_1448), .A2(net_1447), .A1(net_588) );
NOR2_X2 inst_385 ( .A1(net_1434), .A2(net_1062), .ZN(net_916) );
CLKBUF_X2 inst_3319 ( .A(net_2928), .Z(net_3277) );
NOR3_X4 inst_197 ( .A2(net_2343), .A3(net_1358), .ZN(net_1266), .A1(net_548) );
DFFR_X1 inst_2653 ( .D(net_1491), .CK(net_3384), .RN(x2480), .Q(x295) );
CLKBUF_X2 inst_2958 ( .A(net_2915), .Z(net_2916) );
INV_X4 inst_1973 ( .A(net_2257), .ZN(net_1217) );
CLKBUF_X2 inst_3089 ( .A(net_3036), .Z(net_3047) );
OAI22_X2 inst_24 ( .A2(net_1859), .B2(net_1653), .ZN(net_730), .A1(net_728), .B1(net_472) );
CLKBUF_X2 inst_3051 ( .A(net_2944), .Z(net_3009) );
NAND2_X2 inst_1122 ( .ZN(net_667), .A2(net_221), .A1(net_217) );
CLKBUF_X2 inst_3324 ( .A(net_3281), .Z(net_3282) );
NAND2_X2 inst_1209 ( .A2(net_2320), .A1(net_616), .ZN(net_614) );
DFFR_X1 inst_2550 ( .D(net_678), .Q(net_74), .CK(net_2812), .RN(x2480) );
NAND2_X2 inst_1560 ( .ZN(net_2123), .A2(net_2122), .A1(net_2121) );
OAI21_X2 inst_150 ( .ZN(net_1588), .B1(net_1587), .A(net_781), .B2(net_28) );
NAND2_X2 inst_1611 ( .ZN(net_2411), .A1(net_1448), .A2(net_180) );
NAND2_X4 inst_887 ( .ZN(net_1857), .A1(net_907), .A2(net_758) );
CLKBUF_X2 inst_2981 ( .A(net_2891), .Z(net_2939) );
NAND2_X2 inst_1669 ( .ZN(net_2694), .A1(net_2441), .A2(net_2426) );
AOI21_X4 inst_2771 ( .A(net_2548), .B2(net_2360), .B1(net_1720), .ZN(net_1594) );
NAND3_X2 inst_596 ( .A2(net_2267), .A3(net_2061), .ZN(net_822), .A1(net_821) );
NAND2_X2 inst_1663 ( .ZN(net_2665), .A1(net_863), .A2(net_488) );
INV_X4 inst_2142 ( .ZN(net_2205), .A(net_2204) );
AOI22_X2 inst_2714 ( .A2(net_2320), .B1(net_1943), .A1(net_1688), .ZN(net_665), .B2(net_664) );
NAND2_X1 inst_1705 ( .A1(net_632), .ZN(net_100), .A2(x2143) );
CLKBUF_X2 inst_3162 ( .A(net_3119), .Z(net_3120) );
OAI21_X4 inst_90 ( .ZN(net_2172), .B2(net_2171), .B1(net_2169), .A(net_2168) );
NAND2_X4 inst_847 ( .A1(net_2213), .ZN(net_1630), .A2(net_313) );
AOI22_X2 inst_2720 ( .B1(net_2519), .B2(net_994), .ZN(net_879), .A2(net_864), .A1(net_539) );
INV_X2 inst_2357 ( .A(net_1648), .ZN(net_1647) );
NAND2_X1 inst_1716 ( .ZN(net_1123), .A1(net_222), .A2(net_204) );
INV_X4 inst_1942 ( .A(net_1825), .ZN(net_126) );
CLKBUF_X2 inst_3253 ( .A(net_3109), .Z(net_3211) );
DFFR_X1 inst_2648 ( .D(net_1522), .CK(net_3411), .RN(x2480), .Q(x309) );
NAND2_X2 inst_1146 ( .ZN(net_176), .A1(net_137), .A2(net_73) );
INV_X8 inst_1801 ( .ZN(net_1934), .A(net_1933) );
NAND3_X2 inst_637 ( .A1(net_2488), .ZN(net_1660), .A2(net_1421), .A3(net_835) );
NAND4_X2 inst_547 ( .ZN(net_2304), .A4(net_2303), .A3(net_2302), .A2(net_2301), .A1(net_2300) );
CLKBUF_X2 inst_3105 ( .A(net_3062), .Z(net_3063) );
NAND2_X4 inst_720 ( .A1(net_592), .ZN(net_173), .A2(net_108) );
NAND2_X4 inst_958 ( .ZN(net_2260), .A1(net_1585), .A2(net_1484) );
INV_X4 inst_1961 ( .A(net_2578), .ZN(net_707) );
INV_X1 inst_2460 ( .A(net_2415), .ZN(net_1065) );
NAND2_X2 inst_1217 ( .A1(net_1585), .A2(net_1478), .ZN(net_1213) );
INV_X1 inst_2457 ( .A(net_669), .ZN(net_668) );
NOR2_X2 inst_368 ( .A2(net_2561), .A1(net_2129), .ZN(net_705) );
NAND2_X4 inst_1010 ( .ZN(net_2547), .A2(net_2352), .A1(net_2349) );
NAND2_X1 inst_1697 ( .A1(net_2326), .A2(net_1448), .ZN(net_226) );
NAND2_X1 inst_1702 ( .A1(net_1586), .ZN(net_141), .A2(x1889) );
NOR2_X4 inst_274 ( .ZN(net_1751), .A2(net_1750), .A1(net_977) );
NAND2_X2 inst_1277 ( .ZN(net_826), .A1(net_825), .A2(net_585) );
NAND2_X2 inst_1607 ( .ZN(net_2368), .A1(net_2262), .A2(net_2133) );
AOI21_X2 inst_2817 ( .B2(net_2486), .ZN(net_2475), .B1(net_2469), .A(net_1421) );
INV_X4 inst_2092 ( .ZN(net_1719), .A(net_1716) );
NAND2_X4 inst_867 ( .A1(net_1949), .A2(net_1948), .ZN(net_1737) );
OAI21_X2 inst_164 ( .ZN(net_2144), .B1(net_2143), .B2(net_878), .A(net_306) );
CLKBUF_X2 inst_3207 ( .A(net_3164), .Z(net_3165) );
CLKBUF_X2 inst_3027 ( .A(net_2885), .Z(net_2985) );
NAND2_X4 inst_820 ( .ZN(net_1401), .A2(net_1400), .A1(net_976) );
CLKBUF_X2 inst_3143 ( .A(net_3059), .Z(net_3101) );
INV_X4 inst_1854 ( .A(net_1434), .ZN(net_511) );
AOI22_X4 inst_2696 ( .ZN(net_1939), .B2(net_856), .A1(net_243), .A2(net_221), .B1(net_180) );
OAI21_X2 inst_157 ( .A(net_2251), .ZN(net_1854), .B2(net_728), .B1(net_467) );
NAND2_X2 inst_1441 ( .ZN(net_1447), .A1(net_1258), .A2(x1073) );
NAND2_X1 inst_1710 ( .ZN(net_739), .A1(net_736), .A2(net_200) );
CLKBUF_X2 inst_2929 ( .A(net_2886), .Z(net_2887) );
CLKBUF_X2 inst_3443 ( .A(net_3400), .Z(net_3401) );
INV_X2 inst_2407 ( .ZN(net_2701), .A(net_310) );
CLKBUF_X2 inst_2880 ( .A(net_2837), .Z(net_2838) );
INV_X8 inst_1771 ( .A(net_2061), .ZN(net_1158) );
NAND2_X2 inst_1440 ( .A2(net_1686), .ZN(net_1446), .A1(net_1445) );
OAI21_X4 inst_68 ( .B1(net_2568), .B2(net_2169), .ZN(net_1251), .A(net_1026) );
DFFR_X1 inst_2660 ( .D(net_1467), .CK(net_3407), .RN(x2480), .Q(x355) );
CLKBUF_X2 inst_3142 ( .A(net_2883), .Z(net_3100) );
INV_X2 inst_2305 ( .ZN(net_729), .A(net_728) );
INV_X4 inst_1966 ( .ZN(net_2437), .A(net_425) );
CLKBUF_X2 inst_3355 ( .A(net_3312), .Z(net_3313) );
NAND2_X2 inst_1253 ( .ZN(net_725), .A1(net_721), .A2(net_246) );
NAND2_X4 inst_753 ( .A1(net_1229), .A2(net_1025), .ZN(net_758) );
INV_X2 inst_2389 ( .ZN(net_2250), .A(net_2248) );
INV_X4 inst_2150 ( .ZN(net_2297), .A(net_2296) );
CLKBUF_X2 inst_3427 ( .A(net_2938), .Z(net_3385) );
INV_X4 inst_2177 ( .ZN(net_2526), .A(net_2525) );
AOI21_X2 inst_2793 ( .B2(net_1156), .B1(net_899), .ZN(net_834), .A(net_445) );
INV_X4 inst_1884 ( .A(net_2021), .ZN(net_366) );
INV_X4 inst_2018 ( .A(net_2117), .ZN(net_1037) );
INV_X16 inst_2435 ( .ZN(net_2362), .A(net_2361) );
NAND2_X4 inst_946 ( .A2(net_2270), .ZN(net_2189), .A1(net_1084) );
INV_X2 inst_2260 ( .ZN(net_67), .A(x1186) );
INV_X4 inst_1954 ( .A(net_1585), .ZN(net_633) );
INV_X4 inst_2148 ( .ZN(net_2285), .A(net_2284) );
NAND2_X2 inst_1643 ( .A2(net_2587), .ZN(net_2578), .A1(net_769) );
CLKBUF_X2 inst_3410 ( .A(net_3237), .Z(net_3368) );
CLKBUF_X2 inst_2900 ( .A(net_2812), .Z(net_2858) );
NAND2_X1 inst_1690 ( .A2(net_1643), .A1(net_1194), .ZN(net_410) );
INV_X4 inst_2120 ( .ZN(net_1980), .A(net_1978) );
NAND2_X2 inst_1591 ( .A1(net_2587), .ZN(net_2272), .A2(net_1086) );
CLKBUF_X2 inst_3247 ( .A(net_3204), .Z(net_3205) );
NAND2_X2 inst_1678 ( .ZN(net_2719), .A1(net_2718), .A2(net_276) );
NOR2_X2 inst_379 ( .A2(net_1193), .ZN(net_819), .A1(net_818) );
NAND2_X4 inst_926 ( .ZN(net_2083), .A1(net_747), .A2(net_211) );
DFFR_X1 inst_2613 ( .Q(net_2778), .D(net_330), .CK(net_3340), .RN(x2480) );
INV_X4 inst_2053 ( .ZN(net_1297), .A(net_1291) );
OAI22_X4 inst_17 ( .A2(net_2791), .ZN(net_1136), .A1(net_632), .B1(net_133), .B2(net_59) );
NAND2_X2 inst_1325 ( .A1(net_1167), .ZN(net_974), .A2(net_865) );
DFFR_X1 inst_2570 ( .D(net_2760), .CK(net_3271), .RN(x2480), .Q(x159) );
NOR2_X4 inst_249 ( .A2(net_2746), .ZN(net_1230), .A1(net_1227) );
NAND2_X2 inst_1287 ( .ZN(net_1898), .A1(net_86), .A2(x1110) );
INV_X2 inst_2233 ( .ZN(net_300), .A(net_299) );
INV_X2 inst_2234 ( .A(net_2305), .ZN(net_298) );
CLKBUF_X2 inst_3312 ( .A(net_3269), .Z(net_3270) );
NAND2_X2 inst_1169 ( .ZN(net_107), .A1(net_98), .A2(x597) );
NAND2_X2 inst_1649 ( .ZN(net_2600), .A2(net_2597), .A1(net_163) );
NAND2_X4 inst_891 ( .A1(net_1929), .ZN(net_1878), .A2(net_1384) );
NAND2_X2 inst_1480 ( .ZN(net_1723), .A2(net_1722), .A1(net_1721) );
OAI21_X4 inst_74 ( .B1(net_2809), .ZN(net_1564), .A(net_1563), .B2(net_86) );
INV_X2 inst_2244 ( .A(net_1877), .ZN(net_171) );
NAND2_X2 inst_1235 ( .ZN(net_659), .A2(net_586), .A1(net_212) );
NOR2_X4 inst_288 ( .A2(net_2741), .ZN(net_2080), .A1(net_1566) );
NOR2_X2 inst_396 ( .A2(net_1223), .ZN(net_1001), .A1(net_451) );
CLKBUF_X2 inst_3382 ( .A(net_3339), .Z(net_3340) );
CLKBUF_X2 inst_3284 ( .A(net_3241), .Z(net_3242) );
CLKBUF_X2 inst_3046 ( .A(net_2929), .Z(net_3004) );
CLKBUF_X2 inst_3377 ( .A(net_3254), .Z(net_3335) );
CLKBUF_X2 inst_2877 ( .A(net_2834), .Z(net_2835) );
NAND3_X2 inst_669 ( .A2(net_2747), .ZN(net_2233), .A1(net_2232), .A3(net_928) );
NAND3_X2 inst_664 ( .ZN(net_2191), .A1(net_2189), .A2(net_2157), .A3(net_1159) );
NAND2_X2 inst_1298 ( .ZN(net_895), .A1(net_892), .A2(net_210) );
NAND2_X4 inst_917 ( .ZN(net_2022), .A2(net_2017), .A1(net_2001) );
INV_X8 inst_1743 ( .A(net_2386), .ZN(net_319) );
NOR2_X2 inst_372 ( .A1(net_1318), .A2(net_1021), .ZN(net_778) );
NAND2_X2 inst_1600 ( .ZN(net_2337), .A2(net_1962), .A1(net_1961) );
AND2_X2 inst_2850 ( .ZN(net_2369), .A2(net_2368), .A1(net_2367) );
NOR2_X4 inst_215 ( .ZN(net_329), .A1(net_292), .A2(net_287) );
INV_X4 inst_1918 ( .A(net_235), .ZN(net_232) );
AND2_X2 inst_2845 ( .A1(net_2354), .A2(net_1235), .ZN(net_1128) );
NAND2_X2 inst_1418 ( .A1(net_1909), .A2(net_1905), .ZN(net_1363) );
INV_X8 inst_1740 ( .A(net_2111), .ZN(net_345) );
DFFR_X1 inst_2624 ( .Q(net_2757), .D(net_1958), .CK(net_3302), .RN(x2480) );
CLKBUF_X2 inst_2977 ( .A(net_2934), .Z(net_2935) );
NAND2_X4 inst_849 ( .ZN(net_1658), .A1(net_1657), .A2(net_1310) );
NAND2_X2 inst_1092 ( .A2(net_1083), .A1(net_608), .ZN(net_399) );
INV_X2 inst_2397 ( .ZN(net_2457), .A(net_2455) );
INV_X8 inst_1775 ( .A(net_1949), .ZN(net_1240) );
OR2_X4 inst_3 ( .ZN(net_767), .A1(net_766), .A2(net_614) );
NAND2_X2 inst_1172 ( .A1(net_635), .ZN(net_104), .A2(x972) );
INV_X4 inst_2001 ( .A(net_1277), .ZN(net_942) );
NAND2_X2 inst_1090 ( .A1(net_2695), .A2(net_2118), .ZN(net_404) );
CLKBUF_X2 inst_3060 ( .A(net_2895), .Z(net_3018) );
INV_X2 inst_2372 ( .A(net_1820), .ZN(net_1819) );
DFFR_X1 inst_2575 ( .Q(net_2780), .D(net_1299), .CK(net_3041), .RN(x2480) );
NAND2_X2 inst_1657 ( .ZN(net_2624), .A2(net_2621), .A1(net_2273) );
INV_X8 inst_1844 ( .ZN(net_2525), .A(net_2524) );
NAND3_X4 inst_566 ( .A2(net_1089), .ZN(net_595), .A3(net_594), .A1(net_593) );
NAND2_X2 inst_1399 ( .ZN(net_1307), .A2(net_1306), .A1(net_1304) );
NAND2_X2 inst_1239 ( .ZN(net_664), .A2(net_663), .A1(net_662) );
INV_X4 inst_1913 ( .A(net_2106), .ZN(net_248) );
INV_X4 inst_2077 ( .ZN(net_1615), .A(net_1613) );
INV_X2 inst_2368 ( .ZN(net_1769), .A(net_1768) );
INV_X4 inst_1990 ( .ZN(net_854), .A(net_853) );
CLKBUF_X2 inst_3126 ( .A(net_3007), .Z(net_3084) );
AOI22_X2 inst_2735 ( .A2(net_2756), .ZN(net_2035), .A1(net_284), .B1(net_278), .B2(x2026) );
OAI22_X2 inst_36 ( .B2(net_2807), .A2(net_2806), .ZN(net_2743), .B1(net_1008), .A1(net_658) );
CLKBUF_X2 inst_2934 ( .A(net_2891), .Z(net_2892) );
AOI21_X4 inst_2767 ( .A(net_2522), .B1(net_2508), .ZN(net_1186), .B2(net_378) );
NAND2_X2 inst_1370 ( .ZN(net_1188), .A1(net_723), .A2(net_226) );
DFFR_X2 inst_2512 ( .D(net_1836), .Q(net_1526), .CK(net_2908), .RN(x2480) );
NAND4_X4 inst_503 ( .A1(net_2744), .A3(net_2591), .ZN(net_1802), .A4(net_785), .A2(net_784) );
NOR2_X2 inst_451 ( .ZN(net_1992), .A2(net_1114), .A1(net_356) );
INV_X4 inst_2166 ( .ZN(net_2427), .A(net_2426) );
INV_X2 inst_2333 ( .ZN(net_1094), .A(net_546) );
CLKBUF_X2 inst_3193 ( .A(net_3149), .Z(net_3151) );
INV_X4 inst_1936 ( .A(net_647), .ZN(net_140) );
NAND2_X4 inst_797 ( .A2(net_1821), .ZN(net_1231), .A1(net_421) );
NAND2_X2 inst_1495 ( .A1(net_1943), .ZN(net_1758), .A2(net_647) );
INV_X4 inst_2099 ( .ZN(net_1780), .A(net_1779) );
NAND3_X2 inst_686 ( .ZN(net_2617), .A3(net_2616), .A2(net_2271), .A1(net_1713) );
NAND2_X2 inst_1097 ( .A2(net_2408), .ZN(net_355), .A1(net_344) );
CLKBUF_X2 inst_3067 ( .A(net_3014), .Z(net_3025) );
CLKBUF_X2 inst_3032 ( .A(net_2854), .Z(net_2990) );
CLKBUF_X2 inst_2914 ( .A(net_2871), .Z(net_2872) );
INV_X8 inst_1732 ( .A(net_2603), .ZN(net_382) );
CLKBUF_X2 inst_3294 ( .A(net_3251), .Z(net_3252) );
CLKBUF_X2 inst_2888 ( .A(net_2845), .Z(net_2846) );
AOI22_X2 inst_2741 ( .A2(net_2775), .ZN(net_2344), .A1(net_283), .B1(net_126), .B2(x1318) );
NAND2_X4 inst_967 ( .ZN(net_2319), .A1(net_2181), .A2(net_95) );
INV_X4 inst_2119 ( .ZN(net_1975), .A(net_1974) );
NAND2_X2 inst_1522 ( .ZN(net_1947), .A2(net_1604), .A1(net_313) );
INV_X4 inst_1929 ( .A(net_2325), .ZN(net_163) );
INV_X4 inst_1998 ( .ZN(net_922), .A(net_920) );
CLKBUF_X2 inst_3302 ( .A(net_3259), .Z(net_3260) );
CLKBUF_X2 inst_3391 ( .A(net_3348), .Z(net_3349) );
CLKBUF_X2 inst_2870 ( .A(net_2827), .Z(net_2828) );
NAND3_X2 inst_676 ( .A3(net_2506), .ZN(net_2409), .A2(net_2406), .A1(net_2402) );
CLKBUF_X2 inst_3348 ( .A(net_3305), .Z(net_3306) );
INV_X8 inst_1794 ( .ZN(net_1859), .A(net_1858) );
NAND2_X2 inst_1115 ( .A1(net_645), .ZN(net_236), .A2(net_180) );
NAND2_X2 inst_1227 ( .A1(net_1585), .A2(net_1481), .ZN(net_642) );
INV_X2 inst_2324 ( .ZN(net_947), .A(net_946) );
NAND2_X4 inst_874 ( .ZN(net_1786), .A2(net_1735), .A1(net_202) );
CLKBUF_X2 inst_3069 ( .A(net_2911), .Z(net_3027) );
CLKBUF_X2 inst_2976 ( .A(net_2933), .Z(net_2934) );
NAND2_X4 inst_1021 ( .ZN(net_2610), .A1(net_2609), .A2(net_2369) );
NAND2_X2 inst_1681 ( .ZN(net_2730), .A1(net_2729), .A2(net_1918) );
NAND2_X1 inst_1684 ( .A2(net_2406), .A1(net_1180), .ZN(net_519) );
NAND2_X2 inst_1386 ( .ZN(net_1262), .A2(net_174), .A1(net_166) );
INV_X2 inst_2255 ( .ZN(net_225), .A(net_156) );
NAND2_X2 inst_1652 ( .ZN(net_2607), .A2(net_2102), .A1(net_1861) );
NOR2_X4 inst_217 ( .A2(net_1074), .ZN(net_241), .A1(net_240) );
NAND2_X2 inst_1076 ( .A1(net_2423), .A2(net_2160), .ZN(net_470) );
NAND3_X4 inst_572 ( .ZN(net_1902), .A1(net_1787), .A2(net_1234), .A3(net_603) );
NAND2_X2 inst_1622 ( .ZN(net_2482), .A1(net_2481), .A2(net_2204) );
CLKBUF_X2 inst_3047 ( .A(net_3004), .Z(net_3005) );
NAND2_X2 inst_1101 ( .A2(net_1120), .A1(net_913), .ZN(net_336) );
INV_X8 inst_1735 ( .A(net_2288), .ZN(net_360) );
NOR2_X4 inst_257 ( .A1(net_2485), .ZN(net_1419), .A2(net_836) );
INV_X4 inst_2050 ( .A(net_2602), .ZN(net_1280) );
INV_X4 inst_2000 ( .ZN(net_934), .A(net_933) );
CLKBUF_X2 inst_2950 ( .A(net_2907), .Z(net_2908) );
INV_X2 inst_2213 ( .A(net_1193), .ZN(net_402) );
NOR2_X2 inst_485 ( .ZN(net_2628), .A2(net_2603), .A1(net_1286) );
CLKBUF_X2 inst_2897 ( .A(net_2854), .Z(net_2855) );
DFFR_X2 inst_2529 ( .D(net_1571), .Q(net_1477), .CK(net_2956), .RN(x2480) );
NAND2_X4 inst_861 ( .A2(net_2320), .A1(net_1838), .ZN(net_1696) );
NAND2_X2 inst_1195 ( .A2(net_2239), .A1(net_622), .ZN(net_581) );
NAND3_X2 inst_672 ( .ZN(net_2333), .A3(net_1672), .A1(net_845), .A2(net_407) );
NAND2_X2 inst_1471 ( .A1(net_1838), .ZN(net_1691), .A2(net_234) );
INV_X8 inst_1787 ( .ZN(net_1738), .A(net_1737) );
CLKBUF_X2 inst_2990 ( .A(net_2844), .Z(net_2948) );
NAND2_X2 inst_1189 ( .A1(net_2386), .A2(net_856), .ZN(net_574) );
NAND2_X2 inst_1205 ( .A1(net_2308), .A2(net_1462), .ZN(net_604) );
INV_X2 inst_2360 ( .A(net_2293), .ZN(net_1681) );
NAND2_X2 inst_1283 ( .A1(net_1641), .ZN(net_837), .A2(net_499) );
INV_X1 inst_2451 ( .A(net_2113), .ZN(net_372) );
NAND2_X2 inst_1525 ( .ZN(net_1951), .A2(net_198), .A1(net_187) );
CLKBUF_X2 inst_3230 ( .A(net_3187), .Z(net_3188) );
INV_X2 inst_2248 ( .A(net_1191), .ZN(net_157) );
INV_X1 inst_2453 ( .A(net_164), .ZN(net_149) );
NAND2_X2 inst_1202 ( .A2(net_2149), .A1(net_2148), .ZN(net_597) );
NAND2_X2 inst_1312 ( .A1(net_2306), .A2(net_1338), .ZN(net_943) );
NAND2_X2 inst_1540 ( .ZN(net_2012), .A2(net_2010), .A1(net_375) );
CLKBUF_X2 inst_3281 ( .A(net_2970), .Z(net_3239) );
INV_X2 inst_2227 ( .A(net_1567), .ZN(net_348) );
NAND3_X1 inst_703 ( .ZN(net_2549), .A1(net_2548), .A3(net_2295), .A2(net_1927) );
OAI22_X2 inst_33 ( .A2(net_2505), .ZN(net_2430), .B2(net_2408), .B1(net_1632), .A1(net_1429) );
AOI22_X2 inst_2742 ( .A2(net_2772), .ZN(net_2365), .A1(net_283), .B1(net_126), .B2(x1958) );
NAND2_X2 inst_1660 ( .ZN(net_2645), .A1(net_2644), .A2(net_1403) );
NAND3_X2 inst_660 ( .ZN(net_2086), .A1(net_2085), .A3(net_1763), .A2(net_945) );
DFFR_X2 inst_2490 ( .Q(net_1488), .D(net_322), .CK(net_2919), .RN(x2480) );
INV_X4 inst_2107 ( .ZN(net_1835), .A(net_777) );
DFFR_X1 inst_2546 ( .D(net_812), .Q(net_75), .CK(net_3046), .RN(x2480) );
NAND4_X2 inst_517 ( .ZN(net_1044), .A2(net_1043), .A4(net_1005), .A3(net_1003), .A1(net_1002) );
INV_X2 inst_2346 ( .A(net_1428), .ZN(net_1427) );
NAND2_X2 inst_1576 ( .ZN(net_2192), .A1(net_2189), .A2(net_1158) );
NOR2_X4 inst_232 ( .A1(net_1701), .ZN(net_1028), .A2(net_1026) );
NAND2_X2 inst_1261 ( .A2(net_2133), .ZN(net_740), .A1(net_243) );
CLKBUF_X2 inst_3462 ( .A(net_3419), .Z(net_3420) );
CLKBUF_X2 inst_3419 ( .A(net_3376), .Z(net_3377) );
NAND2_X2 inst_1067 ( .A1(net_1272), .A2(net_690), .ZN(net_490) );
NOR2_X4 inst_310 ( .ZN(net_2375), .A2(net_1242), .A1(net_511) );
INV_X8 inst_1824 ( .ZN(net_2328), .A(net_2327) );
NAND2_X2 inst_1214 ( .A1(net_1585), .A2(net_1520), .ZN(net_626) );
NOR2_X4 inst_253 ( .ZN(net_1340), .A2(net_1208), .A1(net_1095) );
NAND2_X4 inst_971 ( .ZN(net_2345), .A2(net_2299), .A1(net_1623) );
NAND2_X2 inst_1417 ( .A1(net_1858), .A2(net_1672), .ZN(net_1356) );
NAND2_X2 inst_1219 ( .ZN(net_2732), .A1(net_1585), .A2(net_1497) );
NAND3_X2 inst_589 ( .A2(net_2048), .A1(net_2047), .ZN(net_288), .A3(net_192) );
AOI222_X1 inst_2754 ( .B1(net_2386), .C2(net_1076), .C1(net_736), .A1(net_721), .A2(net_629), .B2(net_617), .ZN(net_291) );
NAND2_X4 inst_794 ( .A2(net_1666), .ZN(net_1644), .A1(net_1069) );
CLKBUF_X2 inst_3459 ( .A(net_3416), .Z(net_3417) );
NAND2_X4 inst_1005 ( .ZN(net_2520), .A1(net_2518), .A2(net_1168) );
AOI21_X4 inst_2759 ( .A(net_1821), .B2(net_1723), .B1(net_1174), .ZN(net_556) );
NAND2_X2 inst_1147 ( .A2(net_210), .A1(net_203), .ZN(net_174) );
NAND2_X2 inst_1580 ( .ZN(net_2211), .A2(net_210), .A1(net_173) );
INV_X8 inst_1768 ( .ZN(net_1071), .A(net_1069) );
INV_X8 inst_1842 ( .ZN(net_2517), .A(net_2516) );
NAND3_X2 inst_602 ( .A2(net_1230), .ZN(net_907), .A1(net_757), .A3(net_286) );
OAI21_X4 inst_59 ( .ZN(net_848), .A(net_847), .B1(net_137), .B2(net_67) );
INV_X4 inst_1877 ( .A(net_2728), .ZN(net_395) );
CLKBUF_X2 inst_2917 ( .A(net_2874), .Z(net_2875) );
INV_X2 inst_2367 ( .ZN(net_1761), .A(net_1758) );
OAI21_X2 inst_135 ( .B2(net_1284), .ZN(net_1134), .B1(net_865), .A(net_864) );
INV_X16 inst_2423 ( .ZN(net_2071), .A(net_2068) );
CLKBUF_X2 inst_3335 ( .A(net_3163), .Z(net_3293) );
CLKBUF_X2 inst_3256 ( .A(net_3213), .Z(net_3214) );
INV_X2 inst_2351 ( .A(net_2108), .ZN(net_1556) );
NAND2_X4 inst_996 ( .ZN(net_2465), .A1(net_2464), .A2(net_1429) );
NAND2_X2 inst_1408 ( .ZN(net_1333), .A2(net_1332), .A1(net_862) );
CLKBUF_X2 inst_3073 ( .A(net_3030), .Z(net_3031) );
INV_X4 inst_1865 ( .A(net_2339), .ZN(net_424) );
OAI221_X2 inst_37 ( .ZN(net_332), .B1(net_327), .A(net_289), .C2(net_285), .C1(net_170), .B2(net_148) );
INV_X4 inst_1980 ( .ZN(net_811), .A(net_810) );
INV_X4 inst_1853 ( .A(net_1114), .ZN(net_522) );
NAND2_X2 inst_1527 ( .ZN(net_1973), .A2(net_1972), .A1(net_1971) );
INV_X4 inst_1889 ( .A(net_2020), .ZN(net_407) );
NAND2_X2 inst_1664 ( .ZN(net_2671), .A1(net_2667), .A2(net_1509) );
INV_X4 inst_2011 ( .ZN(net_1009), .A(net_1008) );
NAND2_X4 inst_740 ( .A1(net_1585), .A2(net_1523), .ZN(net_662) );
INV_X8 inst_1761 ( .A(net_1008), .ZN(net_721) );
NOR2_X4 inst_264 ( .ZN(net_1460), .A2(net_1420), .A1(net_1419) );
NAND2_X2 inst_1447 ( .ZN(net_1553), .A1(net_1376), .A2(net_239) );
CLKBUF_X2 inst_3117 ( .A(net_2854), .Z(net_3075) );
CLKBUF_X2 inst_2885 ( .A(net_2842), .Z(net_2843) );
DFFR_X1 inst_2632 ( .D(net_69), .CK(net_3362), .RN(x2480), .Q(x223) );
INV_X2 inst_2221 ( .A(net_1724), .ZN(net_368) );
OAI21_X4 inst_84 ( .ZN(net_2042), .B1(net_1083), .B2(net_707), .A(net_607) );
INV_X4 inst_2082 ( .A(net_1652), .ZN(net_1651) );
NAND2_X2 inst_1333 ( .A2(net_1440), .ZN(net_998), .A1(net_403) );
OAI21_X2 inst_173 ( .ZN(net_2508), .B2(net_2507), .A(net_2433), .B1(net_1972) );
INV_X4 inst_1937 ( .A(net_643), .ZN(net_164) );
CLKBUF_X2 inst_3286 ( .A(net_3243), .Z(net_3244) );
AOI22_X2 inst_2709 ( .A2(net_2752), .A1(net_284), .ZN(net_282), .B1(net_278), .B2(x1554) );
NAND3_X2 inst_611 ( .A1(net_2191), .ZN(net_1162), .A3(net_1161), .A2(net_1160) );
NOR2_X4 inst_224 ( .A1(net_1858), .A2(net_1672), .ZN(net_816) );
DFFR_X2 inst_2487 ( .Q(net_1532), .D(net_324), .CK(net_3126), .RN(x2480) );
NAND2_X2 inst_1551 ( .ZN(net_2093), .A1(net_1933), .A2(net_1851) );
CLKBUF_X2 inst_3075 ( .A(net_3032), .Z(net_3033) );
NAND2_X2 inst_1260 ( .ZN(net_738), .A2(net_736), .A1(net_621) );
AOI21_X2 inst_2800 ( .A(net_2165), .ZN(net_1107), .B2(net_703), .B1(net_477) );
NAND2_X2 inst_1088 ( .A2(net_1287), .A1(net_994), .ZN(net_409) );
INV_X2 inst_2406 ( .ZN(net_2677), .A(net_2676) );
NAND2_X4 inst_766 ( .A2(net_2360), .A1(net_1865), .ZN(net_946) );
INV_X4 inst_1943 ( .A(net_633), .ZN(net_143) );
CLKBUF_X2 inst_3270 ( .A(net_3227), .Z(net_3228) );
INV_X4 inst_1908 ( .ZN(net_286), .A(net_270) );
NOR2_X1 inst_490 ( .A1(net_2740), .ZN(net_388), .A2(net_358) );
CLKBUF_X2 inst_3332 ( .A(net_3289), .Z(net_3290) );
CLKBUF_X2 inst_3273 ( .A(net_3230), .Z(net_3231) );
NAND2_X4 inst_801 ( .A2(net_1961), .A1(net_1632), .ZN(net_1248) );
NAND3_X2 inst_692 ( .ZN(net_2679), .A3(net_2676), .A2(net_2674), .A1(net_2673) );
AOI22_X2 inst_2717 ( .A2(net_2757), .ZN(net_842), .A1(net_279), .B1(net_278), .B2(x2211) );
INV_X2 inst_2218 ( .A(net_2740), .ZN(net_442) );
NAND2_X2 inst_1517 ( .A1(net_2516), .A2(net_2407), .ZN(net_1889) );
OAI21_X4 inst_70 ( .B1(net_2373), .A(net_2168), .B2(net_2097), .ZN(net_1257) );
NAND2_X4 inst_870 ( .ZN(net_1750), .A2(net_1238), .A1(net_1237) );
OAI21_X2 inst_129 ( .ZN(net_1019), .A(net_1018), .B2(net_1017), .B1(net_558) );
AOI22_X2 inst_2740 ( .A2(net_2773), .ZN(net_2329), .A1(net_283), .B1(net_126), .B2(x2116) );
NAND2_X2 inst_1309 ( .A1(net_2235), .A2(net_2233), .ZN(net_930) );
NAND2_X2 inst_1531 ( .A2(net_2585), .A1(net_2267), .ZN(net_1984) );
INV_X8 inst_1754 ( .A(net_2132), .ZN(net_585) );
OR2_X2 inst_11 ( .A2(net_2793), .A1(net_1258), .ZN(net_1023) );
CLKBUF_X2 inst_2931 ( .A(net_2888), .Z(net_2889) );
OAI211_X2 inst_188 ( .C2(net_2099), .C1(net_1701), .ZN(net_1574), .B(net_1573), .A(net_1572) );
NAND2_X2 inst_1619 ( .ZN(net_2461), .A2(net_2392), .A1(net_1815) );
CLKBUF_X2 inst_3110 ( .A(net_3067), .Z(net_3068) );
NOR2_X2 inst_441 ( .A2(net_1906), .ZN(net_1668), .A1(net_394) );
CLKBUF_X2 inst_3011 ( .A(net_2968), .Z(net_2969) );
CLKBUF_X2 inst_2922 ( .A(net_2879), .Z(net_2880) );
AOI22_X2 inst_2727 ( .B2(net_2320), .ZN(net_1449), .A2(net_1448), .B1(net_892), .A1(net_721) );
DFFR_X2 inst_2530 ( .Q(net_1531), .D(net_1103), .CK(net_3003), .RN(x2480) );
INV_X2 inst_2276 ( .ZN(net_51), .A(x1636) );
CLKBUF_X2 inst_3183 ( .A(net_3140), .Z(net_3141) );
NAND2_X2 inst_1503 ( .ZN(net_1839), .A2(net_1689), .A1(net_212) );
AND2_X2 inst_2848 ( .ZN(net_1397), .A1(net_1052), .A2(net_281) );
INV_X2 inst_2301 ( .A(net_1021), .ZN(net_570) );
NAND2_X4 inst_808 ( .A2(net_1323), .ZN(net_1291), .A1(net_404) );
NAND2_X2 inst_1537 ( .ZN(net_2003), .A1(net_2002), .A2(x1662) );
NAND2_X4 inst_777 ( .ZN(net_1051), .A1(net_1050), .A2(net_101) );
NAND4_X2 inst_557 ( .ZN(net_2654), .A2(net_2653), .A1(net_2648), .A4(net_1839), .A3(net_1054) );
INV_X4 inst_2041 ( .A(net_2746), .ZN(net_1226) );
NAND2_X4 inst_1037 ( .ZN(net_2721), .A2(net_2130), .A1(net_887) );
NAND2_X2 inst_1383 ( .ZN(net_1894), .A2(net_1250), .A1(net_1249) );
CLKBUF_X2 inst_3279 ( .A(net_3236), .Z(net_3237) );
NAND2_X4 inst_823 ( .A1(net_1585), .A2(net_1504), .ZN(net_1409) );
NAND2_X2 inst_1461 ( .A1(net_1774), .ZN(net_1625), .A2(net_830) );
AND2_X4 inst_2838 ( .ZN(net_2424), .A2(net_1712), .A1(net_1711) );
NAND2_X4 inst_933 ( .ZN(net_2119), .A1(net_1808), .A2(net_1805) );
CLKBUF_X2 inst_3423 ( .A(net_3380), .Z(net_3381) );
CLKBUF_X2 inst_3176 ( .A(net_3133), .Z(net_3134) );
AND2_X4 inst_2833 ( .ZN(net_1893), .A2(net_1738), .A1(net_418) );
NOR2_X4 inst_300 ( .ZN(net_2247), .A1(net_2246), .A2(net_1424) );
NAND2_X2 inst_1250 ( .A2(net_2524), .ZN(net_720), .A1(net_716) );
INV_X4 inst_2042 ( .ZN(net_1227), .A(net_909) );
NAND2_X2 inst_1226 ( .A1(net_1585), .A2(net_1537), .ZN(net_641) );
CLKBUF_X2 inst_3325 ( .A(net_3282), .Z(net_3283) );
NAND2_X4 inst_1013 ( .ZN(net_2560), .A1(net_2460), .A2(net_2101) );
NOR2_X2 inst_446 ( .A2(net_2069), .ZN(net_1799), .A1(net_833) );
NOR2_X2 inst_364 ( .A1(net_1492), .ZN(net_151), .A2(net_146) );
INV_X4 inst_1979 ( .A(net_1407), .ZN(net_807) );
INV_X2 inst_2354 ( .A(net_2517), .ZN(net_1601) );
NOR3_X4 inst_195 ( .ZN(net_797), .A2(net_796), .A3(net_541), .A1(net_474) );
CLKBUF_X2 inst_2997 ( .A(net_2954), .Z(net_2955) );
NAND2_X4 inst_824 ( .A2(net_1927), .A1(net_1452), .ZN(net_1411) );
NOR2_X2 inst_411 ( .A2(net_1298), .ZN(net_1197), .A1(net_1155) );
INV_X4 inst_1987 ( .ZN(net_843), .A(net_842) );
AOI21_X2 inst_2796 ( .B1(net_1164), .ZN(net_985), .B2(net_981), .A(net_363) );
OAI21_X2 inst_124 ( .B2(net_1008), .ZN(net_844), .A(net_196), .B1(net_138) );
NAND2_X2 inst_1150 ( .A1(net_617), .A2(net_180), .ZN(net_162) );
AOI22_X2 inst_2729 ( .B2(net_2328), .A2(net_2133), .B1(net_2030), .ZN(net_1570), .A1(net_244) );
NAND2_X2 inst_1413 ( .ZN(net_1345), .A1(net_1344), .A2(net_309) );
INV_X8 inst_1815 ( .ZN(net_2176), .A(net_2175) );
CLKBUF_X2 inst_3430 ( .A(net_3387), .Z(net_3388) );
NAND2_X2 inst_1270 ( .A1(net_1260), .ZN(net_775), .A2(net_163) );
NAND2_X2 inst_1589 ( .A2(net_2326), .ZN(net_2266), .A1(net_2262) );
CLKBUF_X2 inst_3448 ( .A(net_3405), .Z(net_3406) );
INV_X4 inst_2169 ( .ZN(net_2446), .A(net_2445) );
NAND2_X2 inst_1326 ( .A1(net_2738), .A2(net_1361), .ZN(net_978) );
CLKBUF_X2 inst_3439 ( .A(net_3396), .Z(net_3397) );
OAI21_X4 inst_61 ( .B1(net_1585), .ZN(net_892), .A(net_128), .B2(net_42) );
NOR3_X2 inst_203 ( .A1(net_2268), .A3(net_2164), .ZN(net_1182), .A2(net_1085) );
NAND2_X2 inst_1139 ( .A1(net_2328), .A2(net_825), .ZN(net_190) );
NOR2_X2 inst_335 ( .ZN(net_554), .A1(net_542), .A2(net_524) );
NAND2_X2 inst_1519 ( .A2(net_2237), .ZN(net_1940), .A1(net_1260) );
INV_X4 inst_2156 ( .ZN(net_2352), .A(net_2351) );
DFFR_X1 inst_2629 ( .Q(net_2771), .D(net_928), .CK(net_3089), .RN(x2480) );
NAND2_X2 inst_1571 ( .A2(net_2290), .ZN(net_2166), .A1(net_960) );
NAND3_X2 inst_658 ( .ZN(net_2038), .A2(net_520), .A1(net_470), .A3(net_452) );
DFFR_X2 inst_2515 ( .D(net_2675), .Q(net_1537), .CK(net_2984), .RN(x2480) );
NAND2_X4 inst_832 ( .ZN(net_1548), .A1(net_1547), .A2(net_1021) );
NOR2_X2 inst_456 ( .ZN(net_2032), .A1(net_2031), .A2(net_240) );
NAND2_X2 inst_1402 ( .ZN(net_1314), .A2(net_794), .A1(net_491) );
NAND2_X2 inst_1491 ( .A1(net_2494), .ZN(net_1760), .A2(net_1759) );
NOR2_X4 inst_275 ( .A1(net_2472), .A2(net_2391), .ZN(net_1771) );
OAI21_X2 inst_117 ( .B1(net_2259), .A(net_627), .ZN(net_185), .B2(net_52) );
NOR2_X2 inst_438 ( .A1(net_2219), .ZN(net_1619), .A2(net_1611) );
CLKBUF_X2 inst_3106 ( .A(net_3063), .Z(net_3064) );
NAND2_X2 inst_1341 ( .A1(net_2272), .ZN(net_1047), .A2(net_822) );
INV_X4 inst_2154 ( .ZN(net_2347), .A(net_2346) );
NAND3_X2 inst_587 ( .A3(net_739), .A2(net_580), .ZN(net_292), .A1(net_264) );
NAND3_X2 inst_666 ( .ZN(net_2221), .A3(net_2220), .A1(net_1783), .A2(net_1663) );
OAI21_X2 inst_154 ( .ZN(net_1745), .A(net_872), .B1(net_534), .B2(net_507) );
INV_X16 inst_2416 ( .A(net_1585), .ZN(net_1258) );
DFFR_X1 inst_2602 ( .Q(net_2764), .D(net_2226), .CK(net_2988), .RN(x2480) );
NOR2_X4 inst_324 ( .ZN(net_2585), .A2(net_2584), .A1(net_2583) );
NOR2_X2 inst_465 ( .A2(net_2374), .A1(net_2206), .ZN(net_2114) );
INV_X8 inst_1829 ( .A(net_2647), .ZN(net_2398) );
INV_X2 inst_2304 ( .A(net_715), .ZN(net_714) );
OAI21_X2 inst_109 ( .A(net_799), .ZN(net_540), .B1(net_457), .B2(net_429) );
NAND2_X2 inst_1182 ( .ZN(net_89), .A1(net_86), .A2(x815) );
DFFR_X2 inst_2503 ( .D(net_2278), .Q(net_1535), .CK(net_2863), .RN(x2480) );
OAI221_X1 inst_43 ( .B1(net_2592), .A(net_1830), .C1(net_1733), .ZN(net_328), .B2(net_327), .C2(net_319) );
INV_X4 inst_2128 ( .ZN(net_2024), .A(net_1870) );
NAND2_X1 inst_1707 ( .A2(net_2061), .A1(net_769), .ZN(net_606) );
NAND2_X2 inst_1444 ( .A2(net_2398), .ZN(net_1549), .A1(net_437) );
INV_X4 inst_2173 ( .ZN(net_2499), .A(net_2418) );
NAND2_X2 inst_1231 ( .A1(net_1585), .A2(net_1475), .ZN(net_649) );
OAI21_X4 inst_94 ( .ZN(net_2238), .B1(net_2236), .A(net_1732), .B2(net_164) );
INV_X8 inst_1790 ( .A(net_1822), .ZN(net_1821) );
NOR2_X2 inst_375 ( .ZN(net_792), .A1(net_791), .A2(net_526) );
CLKBUF_X2 inst_3214 ( .A(net_3171), .Z(net_3172) );
NAND2_X4 inst_904 ( .A2(net_2408), .A1(net_2338), .ZN(net_1963) );
CLKBUF_X2 inst_3315 ( .A(net_3272), .Z(net_3273) );
INV_X4 inst_1905 ( .ZN(net_326), .A(net_312) );
INV_X2 inst_2264 ( .ZN(net_63), .A(x1456) );
INV_X4 inst_2159 ( .ZN(net_2384), .A(net_2383) );
NOR2_X4 inst_243 ( .A2(net_1225), .ZN(net_1171), .A1(net_1170) );
NAND2_X2 inst_1378 ( .A1(net_2520), .A2(net_2467), .ZN(net_1220) );
NOR2_X4 inst_285 ( .ZN(net_2021), .A2(net_2017), .A1(net_1652) );
AOI22_X4 inst_2697 ( .ZN(net_2432), .B2(net_1125), .B1(net_1124), .A2(net_1121), .A1(net_1118) );
NAND3_X2 inst_591 ( .ZN(net_273), .A2(net_206), .A3(net_201), .A1(net_194) );
NOR2_X2 inst_424 ( .ZN(net_1370), .A1(net_778), .A2(net_435) );
INV_X8 inst_1830 ( .ZN(net_2406), .A(net_2405) );
CLKBUF_X2 inst_3166 ( .A(net_3123), .Z(net_3124) );
OAI22_X4 inst_15 ( .B2(net_2799), .B1(net_632), .ZN(net_330), .A1(net_137), .A2(net_65) );
NAND2_X4 inst_757 ( .A2(net_2360), .A1(net_1719), .ZN(net_802) );
NOR2_X2 inst_343 ( .A1(net_2513), .A2(net_717), .ZN(net_425) );
NAND2_X2 inst_1627 ( .ZN(net_2492), .A1(net_2481), .A2(net_1432) );
INV_X2 inst_2237 ( .A(net_1173), .ZN(net_281) );
NAND2_X2 inst_1563 ( .ZN(net_2126), .A2(net_1007), .A1(net_216) );
NAND4_X2 inst_543 ( .ZN(net_2039), .A2(net_2026), .A1(net_954), .A4(net_953), .A3(net_447) );
NAND2_X2 inst_1106 ( .A2(net_727), .A1(net_576), .ZN(net_270) );
CLKBUF_X2 inst_3242 ( .A(net_3199), .Z(net_3200) );
CLKBUF_X2 inst_3138 ( .A(net_3095), .Z(net_3096) );
NAND2_X4 inst_982 ( .ZN(net_2382), .A2(net_134), .A1(net_122) );
NAND2_X4 inst_929 ( .A2(net_2561), .ZN(net_2095), .A1(net_2094) );
INV_X4 inst_2070 ( .ZN(net_1560), .A(net_535) );
NAND2_X2 inst_1397 ( .ZN(net_1299), .A2(net_176), .A1(net_141) );
NAND2_X2 inst_1256 ( .A1(net_1585), .A2(net_1477), .ZN(net_732) );
CLKBUF_X2 inst_2890 ( .A(net_2813), .Z(net_2848) );
INV_X4 inst_2123 ( .A(net_2177), .ZN(net_2001) );
NOR2_X4 inst_299 ( .ZN(net_2204), .A2(net_1949), .A1(net_1948) );
CLKBUF_X2 inst_3229 ( .A(net_3062), .Z(net_3187) );
AOI22_X2 inst_2706 ( .A2(net_2767), .ZN(net_306), .B1(net_296), .A1(net_284), .B2(x1343) );
INV_X8 inst_1798 ( .A(net_1908), .ZN(net_1907) );
CLKBUF_X2 inst_2927 ( .A(net_2884), .Z(net_2885) );
NOR2_X2 inst_476 ( .ZN(net_2521), .A2(net_2518), .A1(net_450) );
AND2_X4 inst_2827 ( .ZN(net_1418), .A2(net_1195), .A1(net_1109) );
DFFR_X2 inst_2499 ( .D(net_2195), .Q(net_1533), .CK(net_3232), .RN(x2480) );
CLKBUF_X2 inst_3303 ( .A(net_3260), .Z(net_3261) );
INV_X1 inst_2448 ( .A(net_717), .ZN(net_389) );
OAI22_X4 inst_20 ( .A2(net_2785), .ZN(net_2379), .A1(net_634), .B1(net_143), .B2(net_43) );
NAND2_X2 inst_1369 ( .A1(net_1904), .A2(net_1863), .ZN(net_1176) );
INV_X4 inst_1903 ( .A(net_2105), .ZN(net_333) );
NOR2_X2 inst_349 ( .A2(net_2399), .ZN(net_393), .A1(net_354) );
AOI21_X4 inst_2760 ( .A(net_1356), .B1(net_1080), .ZN(net_541), .B2(net_527) );
DFFR_X1 inst_2541 ( .Q(net_869), .D(net_563), .CK(net_3084), .RN(x2480) );
INV_X4 inst_1938 ( .A(net_587), .ZN(net_136) );
NAND3_X4 inst_576 ( .ZN(net_2213), .A1(net_2212), .A2(net_1781), .A3(net_1780) );
DFFR_X1 inst_2554 ( .QN(net_2785), .Q(net_1491), .D(net_1369), .CK(net_3102), .RN(x2480) );
NAND2_X1 inst_1693 ( .A2(net_1689), .A1(net_631), .ZN(net_265) );
AOI22_X2 inst_2745 ( .A2(net_2766), .ZN(net_2416), .A1(net_295), .B1(net_126), .B2(x1222) );
INV_X4 inst_2095 ( .ZN(net_1733), .A(net_1731) );
CLKBUF_X2 inst_3306 ( .A(net_3263), .Z(net_3264) );
DFFR_X1 inst_2561 ( .QN(net_2790), .Q(net_1524), .D(net_560), .CK(net_3050), .RN(x2480) );
NAND2_X4 inst_1020 ( .ZN(net_2611), .A1(net_2610), .A2(net_2435) );
DFFR_X1 inst_2604 ( .Q(net_2767), .D(net_871), .CK(net_3036), .RN(x2480) );
CLKBUF_X2 inst_3055 ( .A(net_3012), .Z(net_3013) );
CLKBUF_X2 inst_2876 ( .A(net_2833), .Z(net_2834) );
NAND2_X2 inst_1244 ( .A2(net_2320), .ZN(net_2149), .A1(net_645) );
CLKBUF_X2 inst_3260 ( .A(net_3217), .Z(net_3218) );
NAND2_X4 inst_976 ( .ZN(net_2361), .A1(net_1926), .A2(net_1013) );
CLKBUF_X2 inst_3248 ( .A(net_3205), .Z(net_3206) );
CLKBUF_X2 inst_3158 ( .A(net_3115), .Z(net_3116) );
INV_X2 inst_2252 ( .A(net_179), .ZN(net_152) );
NAND2_X2 inst_1279 ( .A2(net_2738), .A1(net_984), .ZN(net_828) );
NAND3_X4 inst_582 ( .ZN(net_2651), .A3(net_2650), .A1(net_2648), .A2(net_1054) );
NAND3_X2 inst_683 ( .ZN(net_2550), .A1(net_2545), .A2(net_1927), .A3(net_421) );
NAND2_X2 inst_1096 ( .A2(net_1911), .A1(net_1906), .ZN(net_356) );
CLKBUF_X2 inst_3269 ( .A(net_2944), .Z(net_3227) );
INV_X4 inst_2186 ( .ZN(net_2644), .A(net_2642) );
INV_X4 inst_1944 ( .A(net_634), .ZN(net_133) );
NOR2_X4 inst_210 ( .A2(net_1450), .A1(net_710), .ZN(net_550) );
CLKBUF_X2 inst_3101 ( .A(net_2896), .Z(net_3059) );
INV_X2 inst_2238 ( .A(net_871), .ZN(net_249) );
AOI21_X4 inst_2763 ( .B1(net_2568), .B2(net_2567), .ZN(net_887), .A(net_808) );
INV_X4 inst_2110 ( .ZN(net_1906), .A(net_1905) );
INV_X4 inst_1850 ( .ZN(net_502), .A(net_501) );
CLKBUF_X2 inst_3151 ( .A(net_2877), .Z(net_3109) );
INV_X8 inst_1839 ( .ZN(net_2505), .A(net_2408) );
INV_X4 inst_1950 ( .A(net_1189), .ZN(net_572) );
NAND2_X4 inst_761 ( .A2(net_1898), .A1(net_1897), .ZN(net_856) );
CLKBUF_X2 inst_3414 ( .A(net_3371), .Z(net_3372) );
CLKBUF_X2 inst_3399 ( .A(net_3356), .Z(net_3357) );
AOI21_X2 inst_2803 ( .B2(net_2730), .A(net_2395), .ZN(net_1208), .B1(net_420) );
NAND2_X2 inst_1294 ( .A2(net_2723), .A1(net_2036), .ZN(net_886) );
NAND2_X1 inst_1712 ( .A1(net_1230), .ZN(net_759), .A2(net_286) );
NAND2_X4 inst_725 ( .A2(net_639), .A1(net_564), .ZN(net_217) );
NAND2_X2 inst_1432 ( .A2(net_2640), .A1(net_2638), .ZN(net_1398) );
INV_X4 inst_2057 ( .A(net_1984), .ZN(net_1329) );
CLKBUF_X2 inst_3108 ( .A(net_2944), .Z(net_3066) );
NAND2_X4 inst_747 ( .ZN(net_722), .A2(net_721), .A1(net_621) );
NAND2_X4 inst_843 ( .A2(net_2562), .A1(net_1702), .ZN(net_1607) );
CLKBUF_X2 inst_2853 ( .A(net_2810), .Z(net_2811) );
INV_X8 inst_1779 ( .A(net_1961), .ZN(net_1429) );
CLKBUF_X2 inst_3084 ( .A(net_2985), .Z(net_3042) );
INV_X4 inst_2115 ( .ZN(net_1921), .A(net_1622) );
INV_X2 inst_2259 ( .ZN(net_68), .A(x1024) );
NAND2_X2 inst_1337 ( .ZN(net_1011), .A1(net_119), .A2(net_109) );
CLKBUF_X2 inst_3251 ( .A(net_3208), .Z(net_3209) );
CLKBUF_X2 inst_3096 ( .A(net_3053), .Z(net_3054) );
DFFR_X1 inst_2641 ( .D(net_78), .CK(net_3132), .RN(x2480), .Q(x459) );
INV_X1 inst_2464 ( .A(net_1650), .ZN(net_1649) );
OAI21_X2 inst_112 ( .B2(net_2132), .ZN(net_263), .A(net_183), .B1(net_157) );
NAND2_X1 inst_1728 ( .ZN(net_2187), .A1(net_2077), .A2(net_835) );
CLKBUF_X2 inst_3015 ( .A(net_2972), .Z(net_2973) );
AOI21_X4 inst_2775 ( .B2(net_2153), .ZN(net_2040), .B1(net_2039), .A(net_2038) );
NAND2_X4 inst_916 ( .A2(net_2111), .ZN(net_2020), .A1(net_2017) );
NAND2_X1 inst_1722 ( .A2(net_1947), .A1(net_1946), .ZN(net_1664) );
CLKBUF_X2 inst_3328 ( .A(net_2965), .Z(net_3286) );
NOR2_X4 inst_305 ( .ZN(net_2299), .A2(net_2298), .A1(net_2292) );
NAND2_X2 inst_1638 ( .ZN(net_2574), .A2(net_2573), .A1(net_2571) );
INV_X16 inst_2441 ( .ZN(net_2562), .A(net_2561) );
CLKBUF_X2 inst_3220 ( .A(net_2863), .Z(net_3178) );
NAND2_X2 inst_1111 ( .A1(net_725), .ZN(net_254), .A2(net_228) );
NAND2_X2 inst_1595 ( .ZN(net_2309), .A2(net_2308), .A1(net_2307) );
DFFR_X1 inst_2658 ( .D(net_1468), .CK(net_3410), .RN(x2480), .Q(x323) );
AOI22_X2 inst_2724 ( .A2(net_2750), .ZN(net_1173), .A1(net_295), .B1(net_126), .B2(x1286) );
NAND2_X4 inst_878 ( .A2(net_1920), .ZN(net_1808), .A1(net_1806) );
DFFR_X2 inst_2525 ( .Q(net_1527), .D(net_1301), .CK(net_2975), .RN(x2480) );
CLKBUF_X2 inst_2968 ( .A(net_2925), .Z(net_2926) );
NOR2_X2 inst_480 ( .ZN(net_2543), .A2(net_2540), .A1(net_921) );
INV_X4 inst_1926 ( .ZN(net_284), .A(net_126) );
CLKBUF_X2 inst_2964 ( .A(net_2921), .Z(net_2922) );
INV_X2 inst_2349 ( .ZN(net_1458), .A(net_381) );
CLKBUF_X2 inst_2986 ( .A(net_2943), .Z(net_2944) );
NAND3_X2 inst_646 ( .ZN(net_1887), .A3(net_1882), .A2(net_1059), .A1(net_855) );
NAND4_X1 inst_564 ( .ZN(net_2723), .A3(net_2722), .A2(net_1670), .A1(net_1599), .A4(net_885) );
INV_X2 inst_2206 ( .A(net_2514), .ZN(net_455) );
CLKBUF_X2 inst_3169 ( .A(net_2850), .Z(net_3127) );
AOI21_X2 inst_2792 ( .B1(net_2363), .A(net_1820), .B2(net_1183), .ZN(net_801) );
NAND2_X4 inst_963 ( .A2(net_2727), .ZN(net_2286), .A1(net_779) );
NAND2_X4 inst_739 ( .A1(net_1585), .A2(net_1521), .ZN(net_637) );
NOR2_X2 inst_382 ( .A1(net_2473), .A2(net_1611), .ZN(net_891) );
INV_X2 inst_2329 ( .A(net_2581), .ZN(net_1064) );
NAND2_X4 inst_907 ( .ZN(net_1970), .A2(net_1969), .A1(net_1968) );
NAND2_X4 inst_934 ( .ZN(net_2130), .A2(net_2129), .A1(net_2128) );
OAI21_X4 inst_46 ( .B1(net_2259), .ZN(net_209), .A(net_114), .B2(net_33) );
DFFR_X1 inst_2537 ( .QN(net_2799), .Q(net_1471), .D(net_562), .CK(net_3355), .RN(x2480) );
NAND2_X4 inst_922 ( .ZN(net_2043), .A2(net_2042), .A1(net_2041) );
NAND2_X4 inst_1000 ( .A1(net_2687), .ZN(net_2480), .A2(net_335) );
NAND2_X2 inst_1614 ( .A1(net_2626), .ZN(net_2417), .A2(net_2416) );
NAND2_X2 inst_1126 ( .ZN(net_2148), .A2(net_1007), .A1(net_622) );
NAND2_X2 inst_1502 ( .A2(net_2237), .ZN(net_1831), .A1(net_1828) );
AOI21_X2 inst_2788 ( .B2(net_2499), .A(net_95), .ZN(net_83), .B1(net_82) );
DFFR_X1 inst_2585 ( .D(net_2781), .CK(net_2847), .RN(x2480), .Q(x429) );
NAND2_X4 inst_796 ( .ZN(net_1219), .A2(net_1202), .A1(net_1031) );
INV_X2 inst_2364 ( .A(net_2362), .ZN(net_1722) );
NAND3_X2 inst_633 ( .A1(net_2188), .A3(net_2139), .A2(net_2012), .ZN(net_1598) );
NAND4_X2 inst_524 ( .A3(net_2576), .A4(net_2247), .ZN(net_1276), .A2(net_1207), .A1(net_942) );
INV_X4 inst_1882 ( .A(net_2603), .ZN(net_532) );
OAI21_X4 inst_104 ( .ZN(net_2593), .A(net_1615), .B2(net_1200), .B1(net_602) );
INV_X2 inst_2285 ( .ZN(net_42), .A(x914) );
INV_X2 inst_2331 ( .A(net_1098), .ZN(net_1074) );
NAND2_X2 inst_1049 ( .ZN(net_551), .A1(net_536), .A2(net_364) );
CLKBUF_X2 inst_3344 ( .A(net_3301), .Z(net_3302) );
CLKBUF_X2 inst_3447 ( .A(net_3404), .Z(net_3405) );
OAI21_X2 inst_168 ( .ZN(net_2307), .B2(net_2248), .B1(net_1999), .A(net_934) );
NAND2_X2 inst_1568 ( .ZN(net_2158), .A2(net_2157), .A1(net_2156) );
NAND2_X2 inst_1499 ( .A2(net_1921), .ZN(net_1805), .A1(net_1804) );
INV_X2 inst_2377 ( .A(net_1904), .ZN(net_1903) );
CLKBUF_X2 inst_2972 ( .A(net_2825), .Z(net_2930) );
DFFR_X2 inst_2522 ( .D(net_1675), .Q(net_1464), .CK(net_2882), .RN(x2480) );
CLKBUF_X2 inst_3366 ( .A(net_3323), .Z(net_3324) );
NAND2_X4 inst_873 ( .ZN(net_1766), .A1(net_1154), .A2(net_510) );
NAND2_X4 inst_727 ( .A1(net_1589), .ZN(net_134), .A2(x1170) );
NAND2_X4 inst_991 ( .ZN(net_2445), .A2(net_1049), .A1(net_797) );
NAND3_X2 inst_653 ( .A1(net_2431), .A2(net_2223), .A3(net_1973), .ZN(net_1965) );
NAND2_X4 inst_882 ( .ZN(net_1838), .A1(net_1837), .A2(net_104) );
CLKBUF_X2 inst_2874 ( .A(net_2831), .Z(net_2832) );
CLKBUF_X2 inst_3297 ( .A(net_3254), .Z(net_3255) );
INV_X16 inst_2431 ( .ZN(net_2323), .A(net_2322) );
NAND3_X4 inst_580 ( .ZN(net_2290), .A2(net_2137), .A1(net_1647), .A3(net_1021) );
OAI21_X2 inst_170 ( .ZN(net_2310), .A(net_1417), .B1(net_517), .B2(net_503) );
INV_X8 inst_1746 ( .A(net_2325), .ZN(net_158) );
CLKBUF_X2 inst_2938 ( .A(net_2895), .Z(net_2896) );
CLKBUF_X2 inst_3371 ( .A(net_3328), .Z(net_3329) );
CLKBUF_X2 inst_3052 ( .A(net_2974), .Z(net_3010) );
NAND2_X4 inst_708 ( .A1(net_2439), .A2(net_1650), .ZN(net_508) );
NAND2_X2 inst_1346 ( .A1(net_2483), .ZN(net_1072), .A2(net_1069) );
NAND2_X2 inst_1374 ( .A2(net_1943), .ZN(net_1199), .A1(net_618) );
NAND2_X4 inst_953 ( .A2(net_2747), .ZN(net_2234), .A1(net_2232) );
INV_X4 inst_1857 ( .A(net_2130), .ZN(net_439) );
CLKBUF_X2 inst_2907 ( .A(net_2840), .Z(net_2865) );
DFFR_X2 inst_2510 ( .D(net_1807), .Q(net_1493), .CK(net_3008), .RN(x2480) );
NAND2_X2 inst_1071 ( .A2(net_2548), .A1(net_1904), .ZN(net_478) );
DFFR_X1 inst_2656 ( .D(net_1517), .CK(net_3379), .RN(x2480), .Q(x237) );
CLKBUF_X2 inst_3000 ( .A(net_2878), .Z(net_2958) );
NAND2_X2 inst_1163 ( .ZN(net_116), .A1(net_115), .A2(net_78) );
NOR2_X2 inst_468 ( .A2(net_2268), .ZN(net_2162), .A1(net_1085) );
NAND2_X2 inst_1099 ( .A2(net_2442), .A1(net_1649), .ZN(net_353) );
NAND2_X2 inst_1421 ( .A2(net_2556), .ZN(net_1369), .A1(net_1368) );
NAND2_X2 inst_1604 ( .ZN(net_2363), .A2(net_2362), .A1(net_2360) );
CLKBUF_X2 inst_3239 ( .A(net_3196), .Z(net_3197) );
CLKBUF_X2 inst_3373 ( .A(net_3113), .Z(net_3331) );
INV_X2 inst_2314 ( .ZN(net_815), .A(net_814) );
INV_X4 inst_2190 ( .ZN(net_2666), .A(net_2665) );
NOR2_X2 inst_429 ( .A1(net_1824), .ZN(net_1416), .A2(net_1411) );
AOI22_X4 inst_2692 ( .B2(net_2557), .ZN(net_1670), .A2(net_1056), .A1(net_1055), .B1(net_479) );
NAND2_X2 inst_1599 ( .ZN(net_2339), .A2(net_2338), .A1(net_2336) );
INV_X4 inst_1994 ( .A(net_1757), .ZN(net_866) );
AOI21_X2 inst_2812 ( .B2(net_2520), .A(net_2433), .B1(net_2409), .ZN(net_2029) );
CLKBUF_X2 inst_3197 ( .A(net_3154), .Z(net_3155) );
INV_X4 inst_2162 ( .ZN(net_2415), .A(net_2414) );
OR2_X2 inst_7 ( .A2(net_1427), .A1(net_1288), .ZN(net_378) );
NOR2_X2 inst_392 ( .ZN(net_945), .A2(net_926), .A1(net_165) );
OAI21_X2 inst_120 ( .B2(net_2551), .ZN(net_701), .B1(net_556), .A(net_517) );
NOR2_X4 inst_294 ( .ZN(net_2141), .A2(net_2140), .A1(net_1239) );
CLKBUF_X2 inst_3450 ( .A(net_3381), .Z(net_3408) );
CLKBUF_X2 inst_3467 ( .A(net_3424), .Z(net_3425) );
DFFR_X1 inst_2593 ( .D(net_2775), .CK(net_3198), .RN(x2480), .Q(x72) );
CLKBUF_X2 inst_3064 ( .A(net_2862), .Z(net_3022) );
NAND2_X2 inst_1514 ( .ZN(net_1882), .A1(net_730), .A2(net_493) );
CLKBUF_X2 inst_3384 ( .A(net_3341), .Z(net_3342) );
INV_X2 inst_2272 ( .ZN(net_55), .A(x870) );
NAND2_X2 inst_1083 ( .A2(net_2165), .ZN(net_447), .A1(net_412) );
NAND3_X4 inst_567 ( .A1(net_2015), .A2(net_1855), .ZN(net_1048), .A3(net_824) );
NAND2_X2 inst_1608 ( .A2(net_2399), .A1(net_2393), .ZN(net_2372) );
CLKBUF_X2 inst_3200 ( .A(net_3157), .Z(net_3158) );
NAND2_X4 inst_810 ( .A2(net_2133), .ZN(net_1316), .A1(net_227) );
NOR2_X4 inst_318 ( .ZN(net_2504), .A1(net_2501), .A2(net_684) );
NAND2_X2 inst_1136 ( .A2(net_2326), .A1(net_629), .ZN(net_195) );
INV_X1 inst_2466 ( .ZN(net_1874), .A(net_1873) );
NOR2_X4 inst_230 ( .A2(net_2153), .ZN(net_991), .A1(net_607) );
NAND2_X2 inst_1484 ( .ZN(net_1732), .A2(net_1731), .A1(net_210) );
NAND2_X2 inst_1601 ( .ZN(net_2341), .A2(net_1998), .A1(net_1353) );
CLKBUF_X2 inst_3035 ( .A(net_2992), .Z(net_2993) );
CLKBUF_X2 inst_2899 ( .A(net_2856), .Z(net_2857) );
NAND2_X4 inst_856 ( .ZN(net_1676), .A1(net_1675), .A2(net_782) );
NAND2_X2 inst_1486 ( .A1(net_2323), .ZN(net_1735), .A2(net_1731) );
INV_X2 inst_2281 ( .ZN(net_46), .A(x1361) );
INV_X4 inst_1893 ( .A(net_2129), .ZN(net_371) );

endmodule
